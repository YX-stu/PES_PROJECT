
----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    14:06:37 04/13/2010 
-- Design Name: 
-- Module Name:    input_ctrl - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;



library basic_lib;


entity input_ctrl is
    port(	clk	:	in std_logic;
			reset	:	in std_logic;
			d_in	: 	in std_logic;
			p_out	:	out std_logic);
end input_ctrl;

-- STUDENT CODE HERE


-- STUDENT CODE until HERE
