library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

--! This testbench tests the rgb2hsv component.

--! The testbench passes several RGB pixels as input to rgb2hsv and checks,
--! if the correspopnding output is correct. In case of unexpected output values,
--! an assertion fault is generated.
entity rgb2hsv_tb is
end entity rgb2hsv_tb;

architecture rtl of rgb2hsv_tb is

    type rgb_t is
        record
            r : STD_LOGIC_VECTOR(7 downto 0);
            g : STD_LOGIC_VECTOR(7 downto 0);
            b : STD_LOGIC_VECTOR(7 downto 0);
        end record;
    type rgb_array_t is array(NATURAL range <>) of rgb_t;

    type hsv_t is
        record
            h : STD_LOGIC_VECTOR(8 downto 0);
            s : STD_LOGIC_VECTOR(7 downto 0);
            v : STD_LOGIC_VECTOR(7 downto 0);
        end record;
    type hsv_array_t is array(NATURAL range <>) of hsv_t;

    signal index : INTEGER := 0;
    signal cycle_counter : INTEGER := 0;

    signal input_start : INTEGER := -1;
    signal output_start : INTEGER := -1;

    constant rgb_data : rgb_array_t := (
        ( "11111111", "00000000", "00000000" ),
        ( "00000000", "11111111", "00000000" ),
        ( "00000000", "00000000", "11111111" ),
        ( "11111111", "11111111", "00000000" ),
        ( "11111111", "00000000", "11111111" ),
        ( "00000000", "11111111", "11111111" ),
        ( "01011100", "11110100", "11000100" ),
        ( "11110111", "00101010", "00011110" ),
        ( "11000110", "10110100", "11100101" ),
        ( "01010101", "00101100", "10011111" ),
        ( "00001011", "01101010", "10010111" ),
        ( "10100110", "01100100", "01011001" ),
        ( "00011111", "01001110", "11101111" ),
        ( "01110001", "11101001", "11110110" ),
        ( "00011100", "10110101", "11111100" ),
        ( "01100000", "00111011", "10000011" ),
        ( "01010000", "01101101", "00110101" ),
        ( "01110011", "00101000", "00101000" ),
        ( "01111010", "10000010", "10100010" ),
        ( "00000110", "00111010", "01110000" ),
        ( "10001101", "01101101", "11011000" ),
        ( "01100110", "01111010", "01110010" ),
        ( "10011100", "11011100", "00010110" ),
        ( "11100111", "10101000", "10111010" ),
        ( "10110111", "10010101", "00101101" ),
        ( "10111101", "00110100", "11000110" ),
        ( "11011110", "00011101", "11111010" ),
        ( "00000111", "10100101", "01101101" ),
        ( "01011100", "00101011", "10010101" ),
        ( "11000010", "00101011", "10010011" ),
        ( "00100001", "00010111", "10000111" ),
        ( "10101101", "10001011", "11110000" ),
        ( "11110100", "10111011", "10011111" ),
        ( "00111110", "10110001", "11010110" ),
        ( "10100000", "10000011", "01000101" ),
        ( "00110010", "10000011", "00110110" ),
        ( "01011010", "10100011", "01011011" ),
        ( "01101001", "11001110", "01100000" ),
        ( "00010101", "10101001", "00001000" ),
        ( "00001000", "01100101", "00100110" ),
        ( "10001000", "11100010", "00000000" ),
        ( "00010100", "11000010", "01101001" ),
        ( "00001100", "01010000", "00101101" ),
        ( "00001000", "11010100", "01000111" ),
        ( "10010111", "00100010", "11000001" ),
        ( "00010100", "10111011", "01010101" ),
        ( "10000110", "11101000", "00010101" ),
        ( "00000000", "10011010", "10101111" ),
        ( "11110101", "00000010", "11101011" ),
        ( "11110000", "11010011", "11000101" ),
        ( "11010001", "11110101", "11100010" ),
        ( "01111100", "01000000", "00101101" ),
        ( "11100111", "10101000", "01000011" ),
        ( "11001110", "01001100", "11100001" ),
        ( "10100101", "10111110", "01110000" ),
        ( "11010011", "11110001", "10110100" ),
        ( "01000010", "10000111", "10011110" ),
        ( "10011011", "00001110", "11100100" ),
        ( "10000011", "00110111", "10010111" ),
        ( "01110101", "10010001", "00001010" ),
        ( "01100101", "01101100", "11000000" ),
        ( "01111001", "01100000", "11100111" ),
        ( "01001010", "00101011", "10011110" ),
        ( "01110011", "00011000", "10110010" ),
        ( "01111010", "11001110", "01111001" ),
        ( "01101101", "11100110", "11110010" ),
        ( "00011010", "10101100", "00000010" ),
        ( "01001110", "00110011", "00010110" ),
        ( "11101101", "01010111", "11111110" ),
        ( "01001000", "11011010", "00111111" ),
        ( "01101101", "10111111", "01100111" ),
        ( "00000100", "00011100", "11111000" ),
        ( "00101011", "10101101", "10000101" ),
        ( "11010101", "10001110", "11010001" ),
        ( "01110011", "01000011", "11011110" ),
        ( "01011000", "10111001", "00011010" ),
        ( "10011111", "10000101", "00100011" ),
        ( "01000101", "00100010", "00110101" ),
        ( "10101101", "00100010", "01011001" ),
        ( "01100001", "11110011", "00101011" ),
        ( "11101001", "11101010", "11101001" ),
        ( "11010111", "10000001", "10010110" ),
        ( "11001100", "10111011", "01101010" ),
        ( "01010101", "01011000", "11110101" ),
        ( "01100000", "11001010", "00111100" ),
        ( "11001010", "10100001", "00000110" ),
        ( "11001011", "10001110", "01000011" ),
        ( "10010111", "11110100", "11000100" ),
        ( "11001010", "11000001", "01110100" ),
        ( "10000111", "11111010", "00001011" ),
        ( "01001010", "00101001", "11101010" ),
        ( "11111110", "01101011", "00011001" ),
        ( "01011010", "00101001", "10111000" ),
        ( "00001010", "01000110", "01101000" ),
        ( "00101101", "01010001", "10111100" ),
        ( "01100110", "01011011", "10001111" ),
        ( "11101010", "01100001", "00011000" ),
        ( "10010001", "01111011", "00101101" ),
        ( "01110101", "01110100", "00100100" ),
        ( "01111100", "11110000", "00001101" ),
        ( "01111001", "01011100", "11101011" ),
        ( "10001000", "00000110", "00000001" ),
        ( "01011101", "01001110", "10011011" ),
        ( "11000101", "11001000", "00101101" ),
        ( "11100111", "01101101", "01101011" ),
        ( "10110011", "01001000", "10101110" ),
        ( "10111000", "11011010", "11100010" ),
        ( "11110000", "00001000", "11101011" ),
        ( "11101111", "01010001", "10001110" ),
        ( "10011100", "01010101", "11101101" ),
        ( "10001001", "01111011", "01111110" ),
        ( "01011101", "10111110", "10010000" ),
        ( "01100100", "01111101", "00100110" ),
        ( "00111110", "11101011", "01110010" ),
        ( "11100100", "01101011", "01110100" ),
        ( "11101100", "01111001", "11100001" ),
        ( "10101111", "10101001", "00111011" ),
        ( "11110011", "10110000", "00111011" ),
        ( "00000100", "01100011", "01000110" ),
        ( "00001010", "00100111", "10000011" ),
        ( "10001000", "10011100", "10101000" ),
        ( "10011011", "10110000", "00010100" ),
        ( "10101100", "10001011", "00101101" ),
        ( "11111001", "00101110", "10110001" ),
        ( "11110011", "00111001", "11110100" ),
        ( "00001101", "00010110", "01101110" ),
        ( "11000001", "10100011", "10010111" ),
        ( "01011111", "11001101", "00100001" ),
        ( "01111110", "11001010", "01110010" ),
        ( "11000010", "00101000", "01100001" ),
        ( "00101000", "01110010", "11100011" ),
        ( "00010010", "10110011", "00110011" ),
        ( "10111000", "10001011", "10011011" ),
        ( "10111111", "10001000", "11111110" ),
        ( "11011101", "01101111", "01011011" ),
        ( "00100001", "11100000", "01011011" ),
        ( "11110100", "01111010", "10101010" ),
        ( "11000011", "10101001", "11011001" ),
        ( "01010100", "10101110", "01110001" ),
        ( "00100110", "10111011", "11010000" ),
        ( "00111111", "01011100", "01111001" ),
        ( "10110001", "10001110", "11010110" ),
        ( "00010100", "00001100", "00111101" ),
        ( "11001010", "01110100", "01110101" ),
        ( "10011110", "00010011", "10011011" ),
        ( "00111111", "11001010", "00110011" ),
        ( "10010000", "10011101", "00110111" ),
        ( "10011000", "10011100", "00000111" ),
        ( "10001100", "00011110", "10111001" ),
        ( "11100000", "10110011", "11010110" ),
        ( "01001000", "01010101", "00110000" ),
        ( "00000110", "00000010", "10001000" ),
        ( "10110010", "01110000", "00110001" ),
        ( "11101110", "11101000", "11010111" ),
        ( "00100000", "11110101", "10010110" ),
        ( "11000000", "11010000", "11101011" ),
        ( "11101000", "01110110", "11101100" ),
        ( "00011011", "00000110", "01010000" ),
        ( "11111111", "00111001", "11101000" ),
        ( "00110110", "11100101", "00000000" ),
        ( "01101100", "01100010", "10000000" ),
        ( "00011001", "10100110", "01100100" ),
        ( "10101100", "00111111", "01110111" ),
        ( "01101001", "01110100", "10100001" ),
        ( "01100001", "10111100", "10000110" ),
        ( "10000111", "10011001", "10001101" ),
        ( "11100100", "00111001", "01011110" ),
        ( "11110010", "11011101", "00011101" ),
        ( "10001010", "00101011", "00111100" ),
        ( "00011111", "01100111", "00101010" ),
        ( "10111111", "01010101", "11000011" ),
        ( "01010011", "11001010", "11100011" ),
        ( "01000111", "10000000", "01011101" ),
        ( "00011101", "00000100", "01001000" ),
        ( "01000100", "11101100", "01001111" ),
        ( "10000001", "10001101", "01110011" ),
        ( "11001111", "00000011", "00111111" ),
        ( "11110010", "11010100", "10101111" ),
        ( "01001001", "11101010", "11101010" ),
        ( "10110000", "10111001", "10000010" ),
        ( "10101111", "00000001", "00101110" ),
        ( "00101001", "11100001", "00101111" ),
        ( "10010000", "01111101", "10111011" ),
        ( "01100001", "11111110", "01101011" ),
        ( "10000010", "10010101", "00001000" ),
        ( "10011000", "01011011", "00101100" ),
        ( "00011111", "00000000", "01011111" ),
        ( "10101001", "01001001", "11011110" ),
        ( "11110001", "10110110", "00011010" ),
        ( "11001011", "01001111", "01101000" ),
        ( "11011111", "00101001", "01101000" ),
        ( "11000011", "00011100", "11000010" ),
        ( "11101110", "10000001", "00111001" ),
        ( "10101101", "10101011", "00001111" ),
        ( "01111000", "01110010", "00011000" ),
        ( "11011001", "00101010", "01101101" ),
        ( "00101100", "11000111", "00100011" ),
        ( "01111000", "01110010", "00000111" ),
        ( "01101011", "11000100", "01011110" ),
        ( "00001110", "00110110", "00001000" ),
        ( "11100001", "11011001", "00010110" ),
        ( "11011110", "00111011", "01111001" ),
        ( "01110000", "01101001", "00010001" ),
        ( "11001110", "00101101", "00111100" ),
        ( "10111111", "10010011", "10110001" ),
        ( "01110111", "11101111", "10011010" ),
        ( "00010001", "00110011", "01101011" ),
        ( "01011001", "10000000", "00100001" ),
        ( "00101111", "10100110", "00001011" ),
        ( "01101101", "11000011", "10111111" ),
        ( "10000111", "11101001", "11000111" ),
        ( "10001101", "11000111", "01100111" ),
        ( "11001111", "00101010", "00010010" ),
        ( "01100110", "01110010", "10100000" ),
        ( "11010011", "11110010", "10011110" ),
        ( "11110100", "10010011", "11000101" ),
        ( "00101110", "01100011", "00100101" ),
        ( "10110010", "10111111", "11101011" ),
        ( "00100000", "01000100", "10111111" ),
        ( "00001101", "10010011", "10100010" ),
        ( "11000110", "11010010", "11110011" ),
        ( "10110101", "00101010", "00001100" ),
        ( "01011000", "10001101", "11001110" ),
        ( "11011110", "11101001", "00000001" ),
        ( "00111010", "01111110", "10010101" ),
        ( "10010110", "11110001", "00111010" ),
        ( "00000101", "10100011", "11111110" ),
        ( "10111001", "11001110", "10110010" ),
        ( "11010001", "10000100", "11101010" ),
        ( "00101000", "01001001", "11000100" ),
        ( "01101001", "00101001", "00010010" ),
        ( "01001110", "01100100", "10110110" ),
        ( "00110001", "11011100", "00110011" ),
        ( "00011000", "11011101", "10011101" ),
        ( "11011111", "10000010", "10010001" ),
        ( "11110001", "11011010", "11110010" ),
        ( "01011111", "01101101", "11101110" ),
        ( "01011000", "10000111", "00100110" ),
        ( "01110100", "11111010", "01001000" ),
        ( "00101100", "11000110", "00010111" ),
        ( "11110110", "01010100", "11110111" ),
        ( "11001010", "01001101", "00111011" ),
        ( "11000001", "00110010", "00000101" ),
        ( "10000111", "10111110", "11010000" ),
        ( "10100110", "01110000", "11011011" ),
        ( "00110000", "10011110", "10000000" ),
        ( "00001011", "11001100", "10010001" ),
        ( "10010110", "00111000", "00101101" ),
        ( "11110000", "00110001", "01111111" ),
        ( "01010011", "11001101", "11101011" ),
        ( "10011100", "01010111", "11101110" ),
        ( "01000100", "10100011", "01001111" ),
        ( "00100000", "10100001", "11110010" ),
        ( "01110010", "11001101", "10010101" ),
        ( "01100011", "01111101", "11010001" ),
        ( "01011110", "11000110", "01010101" ),
        ( "10001010", "10110011", "10001110" ),
        ( "11101101", "00101110", "10111101" ),
        ( "11001010", "01101010", "01100010" ),
        ( "01100011", "01010111", "10000101" ),
        ( "00001000", "11001010", "01010100" ),
        ( "00110001", "01011000", "00011100" ),
        ( "11010111", "01111110", "00110010" ),
        ( "10001001", "11011110", "10111110" ),
        ( "10110010", "10001100", "10001001" ),
        ( "11100110", "00000110", "01110000" ),
        ( "10000110", "00110111", "01111100" ),
        ( "00010010", "11001100", "00011101" ),
        ( "11011111", "11101000", "10001100" ),
        ( "01010111", "00000100", "01000010" ),
        ( "01100100", "01011000", "10100000" ),
        ( "11010000", "11010111", "11101101" ),
        ( "01011100", "01100101", "11111010" ),
        ( "00100001", "00101100", "11111010" ),
        ( "01101111", "01011110", "11011100" ),
        ( "11110110", "10010111", "11010100" ),
        ( "11101100", "10101101", "00000100" ),
        ( "00011110", "10011101", "00100110" ),
        ( "00101101", "00100011", "01001100" ),
        ( "00100001", "01100110", "00111011" ),
        ( "11111111", "01011000", "00001111" ),
        ( "10010100", "00111110", "00000110" ),
        ( "00001011", "11010011", "00100100" ),
        ( "10100110", "01110100", "11111110" ),
        ( "10110101", "11111101", "10001100" ),
        ( "10011001", "01110010", "01011010" ),
        ( "11110111", "00001111", "00101011" ),
        ( "00011101", "00101000", "01010100" ),
        ( "00010101", "01110110", "00011010" ),
        ( "11001001", "00011100", "01101111" ),
        ( "01000000", "01100000", "01111010" ),
        ( "00101101", "10111110", "00000000" ),
        ( "10001001", "01110010", "11011001" ),
        ( "00101011", "11010101", "01100111" ),
        ( "10101100", "11011110", "01110110" ),
        ( "10011001", "00011101", "10111000" ),
        ( "10011101", "01000001", "00010000" ),
        ( "01011111", "01101100", "11001000" ),
        ( "11011011", "00100000", "00001011" ),
        ( "10001010", "11111001", "11010101" ),
        ( "11111000", "11011011", "00000010" ),
        ( "00001100", "10011110", "01000111" ),
        ( "11011010", "01100101", "00101010" ),
        ( "00011110", "00101001", "00111100" ),
        ( "10011010", "00110001", "00001100" ),
        ( "10001000", "00010110", "11010110" ),
        ( "00001011", "00000011", "10000100" ),
        ( "00110010", "01001010", "10001100" ),
        ( "01010111", "10110111", "00000011" ),
        ( "11001001", "10100111", "11101011" ),
        ( "00110011", "00010000", "10000111" ),
        ( "01101011", "10010100", "10001000" ),
        ( "10010011", "00110000", "11001100" ),
        ( "10001011", "11001000", "00010010" ),
        ( "11100100", "01001111", "10011001" ),
        ( "10001010", "11111011", "11000110" ),
        ( "00111110", "10111100", "00111100" ),
        ( "11000010", "01010000", "10110101" ),
        ( "00001101", "01011101", "10010011" ),
        ( "11110001", "10001001", "10011000" ),
        ( "00010011", "00100000", "00110001" ),
        ( "01000010", "01110010", "00101001" ),
        ( "11011110", "00011100", "10000000" ),
        ( "01110000", "11111011", "00111010" ),
        ( "00001100", "01010101", "11110000" ),
        ( "10101100", "11111010", "11111101" ),
        ( "11100001", "01011110", "10010110" ),
        ( "01010100", "10011001", "00111101" ),
        ( "00101000", "01010010", "11000001" ),
        ( "10011011", "11001001", "01111110" ),
        ( "01010110", "11010101", "01110100" ),
        ( "10110001", "01011010", "00110011" ),
        ( "01100000", "00011101", "11001001" ),
        ( "00001111", "10001101", "10001101" ),
        ( "11001110", "00111010", "10011101" ),
        ( "11101110", "00110111", "10011011" ),
        ( "11100110", "00001111", "00100111" ),
        ( "00011001", "11000101", "10100101" ),
        ( "00001010", "10111100", "00110101" ),
        ( "10010010", "11001110", "00001110" ),
        ( "10100000", "01100111", "01010001" ),
        ( "11001000", "11110101", "00100111" ),
        ( "00010101", "10101010", "11111010" ),
        ( "01001110", "00111011", "10101011" ),
        ( "11100100", "00010001", "10101111" ),
        ( "01010010", "00100101", "11101000" ),
        ( "10100000", "01100100", "10000101" ),
        ( "01001010", "00110011", "10111111" ),
        ( "01110100", "10110111", "01111000" ),
        ( "10000110", "10011110", "11111100" ),
        ( "10011101", "01111110", "11000001" ),
        ( "10110011", "01100001", "10111000" ),
        ( "10111011", "00001001", "11001100" ),
        ( "01110001", "11101000", "11000100" ),
        ( "00011101", "00110110", "10101010" ),
        ( "10000100", "00000101", "01001100" ),
        ( "01001001", "01001000", "00010010" ),
        ( "01001110", "11111110", "00110101" ),
        ( "01101110", "00011000", "01001010" ),
        ( "10010011", "11001001", "11100100" ),
        ( "10001100", "00011001", "10010100" ),
        ( "10110011", "11010011", "01101010" ),
        ( "01110000", "11101111", "11110001" ),
        ( "11011111", "11100110", "01001110" ),
        ( "11010001", "10000111", "01011000" ),
        ( "11111001", "00001010", "01101100" ),
        ( "00110111", "11101110", "10110011" ),
        ( "00011000", "01110111", "10100010" ),
        ( "01111010", "01011000", "01000000" ),
        ( "11101011", "11110000", "01000000" ),
        ( "11100111", "00011110", "00100111" ),
        ( "01101111", "00011100", "01110100" ),
        ( "01111111", "10010101", "01100101" ),
        ( "10110011", "10111101", "00110010" ),
        ( "11001011", "00001010", "01011101" ),
        ( "10100000", "11010010", "00111100" ),
        ( "00101010", "01010011", "10101111" ),
        ( "00000001", "00001011", "01100000" ),
        ( "10110110", "10101001", "00100000" ),
        ( "00111100", "00010010", "00000010" ),
        ( "00001101", "11000110", "10111000" ),
        ( "01111100", "10010110", "10001000" ),
        ( "10011110", "10001011", "01101101" ),
        ( "00111010", "00100111", "01001101" ),
        ( "01000111", "10001000", "11100010" ),
        ( "01101101", "00110101", "00010110" ),
        ( "01110101", "01000111", "00110010" ),
        ( "11000000", "11010100", "01001100" ),
        ( "11111000", "00100110", "10110111" ),
        ( "10101000", "00011001", "01101000" ),
        ( "01001010", "00100011", "01001010" ),
        ( "00101110", "00100110", "01000101" ),
        ( "00000010", "11101100", "10000000" ),
        ( "10111110", "01000100", "01100100" ),
        ( "10100000", "00000101", "10111000" ),
        ( "01101100", "10010101", "00111110" ),
        ( "00000001", "11110001", "00101000" ),
        ( "01100001", "01001011", "00111100" ),
        ( "00001110", "10011001", "00100011" ),
        ( "01110100", "01100010", "11101010" ),
        ( "10001100", "01100100", "01010010" ),
        ( "00010111", "01001111", "01111111" ),
        ( "00011000", "11000011", "10010010" ),
        ( "00100001", "00101100", "11010110" ),
        ( "10101100", "00011000", "10110111" ),
        ( "00100010", "00111000", "01100011" ),
        ( "01001011", "01000111", "01101000" ),
        ( "00111001", "11010010", "11010011" ),
        ( "10011101", "01001110", "11000101" ),
        ( "10101110", "00110100", "01010001" ),
        ( "10011111", "10110110", "10100010" ),
        ( "10111001", "10010000", "10100110" ),
        ( "11000011", "11000001", "01110101" ),
        ( "00111100", "01101111", "10110001" ),
        ( "00001000", "10011011", "01001111" ),
        ( "01100000", "01010100", "11101110" ),
        ( "11101110", "11110111", "01101101" ),
        ( "01001110", "00010011", "11110111" ),
        ( "01011101", "11100110", "01001111" ),
        ( "01111110", "01100001", "01010100" ),
        ( "11010010", "11000110", "01010110" ),
        ( "01010011", "10000010", "11101110" ),
        ( "01101110", "10010111", "01001111" ),
        ( "11111101", "00100111", "11111001" ),
        ( "11000000", "00100100", "01111110" ),
        ( "11010100", "11010010", "01000011" ),
        ( "01011111", "10101111", "00000011" ),
        ( "10101111", "01100001", "00011100" ),
        ( "10101010", "00110011", "10110000" ),
        ( "11011111", "10001001", "01010100" ),
        ( "01001010", "01010011", "10100101" ),
        ( "11011001", "01101111", "00001010" ),
        ( "01010110", "10001011", "01010010" ),
        ( "10110100", "10011010", "00111010" ),
        ( "00010101", "01000010", "10101110" ),
        ( "00000000", "11110100", "01001011" ),
        ( "11100000", "11001010", "11000001" ),
        ( "10101110", "10011111", "00010011" ),
        ( "10010000", "01111001", "11010100" ),
        ( "11110011", "10110011", "00001001" ),
        ( "01110101", "01011001", "11101001" ),
        ( "01110011", "01010110", "10010100" ),
        ( "11010010", "00100011", "01000011" ),
        ( "00011001", "10100110", "11000011" ),
        ( "01001101", "10000000", "00100111" ),
        ( "01011111", "01100001", "11001111" ),
        ( "11010100", "11000110", "00011111" ),
        ( "11111011", "01100000", "00110011" ),
        ( "11101000", "10101100", "01100010" ),
        ( "00101100", "00111001", "01000001" ),
        ( "01001110", "10101011", "00111000" ),
        ( "00010100", "10100100", "01111100" ),
        ( "10001101", "11111111", "01100111" ),
        ( "11100110", "01110011", "00011111" ),
        ( "11010001", "10001101", "00001111" ),
        ( "11010111", "01000101", "10010111" ),
        ( "00000000", "00011000", "10000101" ),
        ( "00001110", "00110111", "11100000" ),
        ( "00100101", "10000101", "00001001" ),
        ( "00000001", "01000000", "11111111" ),
        ( "10000010", "00100100", "01101001" ),
        ( "00001100", "11111101", "00001101" ),
        ( "11100100", "00110101", "11110001" ),
        ( "00100001", "00010111", "10011010" ),
        ( "00001110", "00100101", "00111011" ),
        ( "11011010", "10001001", "01001000" ),
        ( "01010111", "00110011", "10110100" ),
        ( "01100100", "01101111", "11101011" ),
        ( "11010001", "10000001", "11111000" ),
        ( "11101110", "00101000", "10011011" ),
        ( "10010000", "10111000", "01010111" ),
        ( "10100101", "11101100", "01110101" ),
        ( "11101010", "11001101", "00010010" ),
        ( "01100111", "00101011", "00000010" ),
        ( "11001000", "10001001", "00111011" ),
        ( "10110011", "01001100", "01110010" ),
        ( "01100010", "11011010", "01000101" ),
        ( "01111011", "10100100", "00111010" ),
        ( "11111010", "00100100", "10010101" ),
        ( "11100100", "11000010", "10110100" ),
        ( "01101110", "00000000", "10111011" ),
        ( "00100000", "01011111", "11001010" ),
        ( "10111111", "00101110", "00100111" ),
        ( "11011011", "10010100", "11011010" ),
        ( "11100011", "10101010", "01100011" ),
        ( "11111001", "00100011", "01010010" ),
        ( "01101100", "00011100", "01000011" ),
        ( "10010110", "11110111", "10110111" ),
        ( "11111001", "00100010", "10001110" ),
        ( "10000011", "00101010", "00010011" ),
        ( "01101001", "00100000", "00000010" ),
        ( "10111010", "00101010", "11111111" ),
        ( "01000011", "10011101", "11001011" ),
        ( "01111111", "11011101", "10111111" ),
        ( "11010100", "01010110", "11000000" ),
        ( "00100010", "11010001", "00110011" ),
        ( "11101110", "10001001", "00000011" ),
        ( "10100010", "11010100", "10000010" ),
        ( "01010110", "00101111", "11011010" ),
        ( "10100100", "10010011", "11001110" ),
        ( "00111001", "00010110", "11010111" ),
        ( "01111010", "00001100", "01010001" ),
        ( "01000100", "00011101", "10101011" ),
        ( "00100110", "11110110", "10110000" ),
        ( "00110100", "00000010", "00111000" ),
        ( "10100011", "01101010", "01110001" ),
        ( "11111000", "01111111", "11000011" ),
        ( "11100001", "01111001", "11001010" ),
        ( "10111100", "10101001", "01001000" ),
        ( "00101011", "01110000", "01001001" ),
        ( "01110001", "11001110", "01101001" ),
        ( "11110011", "11110010", "00001010" ),
        ( "10110110", "01001011", "01110000" ),
        ( "01000001", "00111101", "01101100" ),
        ( "00101001", "00001000", "01010011" ),
        ( "00101011", "00101010", "10001000" ),
        ( "10001010", "10011111", "11000010" ),
        ( "00100100", "11001010", "11100001" ),
        ( "00110110", "01011101", "10100100" ),
        ( "00010000", "10110110", "11110010" ),
        ( "11100010", "10011000", "10010000" ),
        ( "01001011", "01100011", "10110100" ),
        ( "10100100", "00010111", "00100110" ),
        ( "00110010", "00011000", "00110101" ),
        ( "10100100", "01110111", "01001101" ),
        ( "11010000", "01100011", "11000010" ),
        ( "00010001", "11001111", "11001000" ),
        ( "10110101", "00010110", "01101100" ),
        ( "00101101", "00010001", "10100010" ),
        ( "00100010", "00110011", "11000001" ),
        ( "10001001", "11001101", "01011001" ),
        ( "00011010", "01011001", "00001101" ),
        ( "11001110", "01100001", "11010100" ),
        ( "11101011", "10000100", "10001101" ),
        ( "10100011", "10111111", "10000110" ),
        ( "01001111", "01001000", "01010001" ),
        ( "10001011", "01010000", "01010101" ),
        ( "00111110", "11001011", "10111010" ),
        ( "11011011", "10011101", "00010001" ),
        ( "11111001", "00100110", "11100011" ),
        ( "00010010", "11000011", "10100111" ),
        ( "00000100", "11111101", "01010101" ),
        ( "00110010", "11011011", "01010011" ),
        ( "00000000", "01101010", "11001100" ),
        ( "11111001", "11100101", "01111001" ),
        ( "10101000", "10001100", "11111101" ),
        ( "00000100", "11010000", "11110100" ),
        ( "01011100", "01011101", "10011110" ),
        ( "00111100", "10110110", "11111011" ),
        ( "00000000", "10100000", "00100010" ),
        ( "00101000", "01100110", "11101000" ),
        ( "00011110", "11111010", "11011111" ),
        ( "11110101", "11010011", "10000100" ),
        ( "01111110", "10011010", "10011011" ),
        ( "01001101", "00000011", "10101101" ),
        ( "11000001", "00000010", "10110111" ),
        ( "01011101", "10001000", "01100111" ),
        ( "10011000", "11000101", "01101110" ),
        ( "10010011", "10110110", "11000010" ),
        ( "10110001", "01011101", "11011101" ),
        ( "00000010", "00010011", "00010010" ),
        ( "01110100", "01011110", "11011010" ),
        ( "01101001", "10100101", "01101010" ),
        ( "00011100", "10111000", "10111111" ),
        ( "01001010", "00111001", "01100111" ),
        ( "11011000", "11000111", "10101001" ),
        ( "10100101", "10110110", "10100010" ),
        ( "11111000", "01011011", "11110000" ),
        ( "00100111", "00001110", "01011110" ),
        ( "01010000", "00000110", "10110100" ),
        ( "11101001", "01111100", "01011111" ),
        ( "01010100", "01001010", "11010101" ),
        ( "00011100", "00000000", "11011011" ),
        ( "10100000", "10000011", "10110110" ),
        ( "00110100", "01100100", "00001011" ),
        ( "11100011", "10011111", "10010010" ),
        ( "01101111", "00100101", "11001101" ),
        ( "01101011", "00000010", "01010101" ),
        ( "11000111", "00011111", "01000010" ),
        ( "11000101", "00100110", "00110010" ),
        ( "10101111", "11000110", "10000111" ),
        ( "00100100", "11011110", "01101110" ),
        ( "00111010", "01010001", "11001001" ),
        ( "10011000", "00111010", "00010110" ),
        ( "01101001", "00101011", "01100010" ),
        ( "00110101", "10000111", "10100000" ),
        ( "11011101", "01111011", "11001111" ),
        ( "10111110", "11011111", "10100000" ),
        ( "00100110", "10101000", "10010010" ),
        ( "01101110", "00111101", "00011010" ),
        ( "01010100", "00100101", "01100110" ),
        ( "11110000", "00011111", "00011111" ),
        ( "10100111", "11101000", "01001000" ),
        ( "10110000", "00001101", "10101000" ),
        ( "01101101", "01010000", "01000011" ),
        ( "00000011", "10101001", "11111100" ),
        ( "01100011", "01111000", "00001001" ),
        ( "11011001", "00001100", "11111011" ),
        ( "01000100", "00011011", "10110101" ),
        ( "11111001", "10100110", "00100101" ),
        ( "01000001", "10010110", "01001110" ),
        ( "11110001", "11010011", "00111001" ),
        ( "10011001", "10110011", "11100011" ),
        ( "01001010", "11011110", "10111001" ),
        ( "10010010", "00111010", "01011100" ),
        ( "10010110", "00111010", "11000100" ),
        ( "01110000", "01111111", "01001010" ),
        ( "01110011", "00001100", "11110101" ),
        ( "01010001", "01100101", "01100100" ),
        ( "10100101", "01011000", "01001110" ),
        ( "11101010", "10001100", "01110101" ),
        ( "10111111", "01111101", "01011110" ),
        ( "10011101", "10101001", "11011101" ),
        ( "00101001", "10111010", "00011101" ),
        ( "01100011", "00110101", "11111101" ),
        ( "01010101", "11101111", "00110000" ),
        ( "01110110", "11111000", "00100001" ),
        ( "10000111", "11100010", "10011010" ),
        ( "11001100", "00010111", "11000100" ),
        ( "10000010", "10100111", "00000101" ),
        ( "10110111", "10110001", "01000110" ),
        ( "11101010", "00000010", "00100000" ),
        ( "01001001", "00110100", "01101101" ),
        ( "01001000", "11010100", "11001001" ),
        ( "01010011", "11100111", "00111111" ),
        ( "11101101", "11111001", "00000010" ),
        ( "00001110", "01100101", "00011110" ),
        ( "00100110", "00100011", "11011100" ),
        ( "11010011", "11110100", "00110010" ),
        ( "10000111", "10001101", "11011101" ),
        ( "01110110", "00000101", "01111001" ),
        ( "00101001", "10100010", "10001001" ),
        ( "00001111", "00111110", "00011011" ),
        ( "00111010", "11101010", "00011111" ),
        ( "01100100", "11011010", "11010111" ),
        ( "00110011", "11011001", "10100110" ),
        ( "00101100", "01001000", "10100001" ),
        ( "01111110", "01011011", "11010111" ),
        ( "11011110", "01000110", "11000110" ),
        ( "10001001", "00100110", "10001100" ),
        ( "11010101", "11111011", "00110111" ),
        ( "01101011", "01000110", "10111110" ),
        ( "11100110", "10101111", "11000101" ),
        ( "10100011", "01011001", "00111001" ),
        ( "10111101", "00110101", "01110110" ),
        ( "10100110", "01101101", "10000110" ),
        ( "10011011", "00101011", "00111110" ),
        ( "00101111", "10010000", "11000011" ),
        ( "01010100", "10010010", "10111010" ),
        ( "10001101", "01100011", "01100010" ),
        ( "10010001", "01101111", "11000100" ),
        ( "01100110", "01010100", "00000000" ),
        ( "11001000", "01111001", "11111011" ),
        ( "10100101", "01001100", "11010110" ),
        ( "01101101", "11111010", "10001101" ),
        ( "10010010", "11110011", "01110011" ),
        ( "00111110", "01101010", "11101100" ),
        ( "01000011", "11011000", "10111111" ),
        ( "11000011", "01111100", "00110010" ),
        ( "11011111", "00011111", "01111000" ),
        ( "01010001", "10000110", "01011001" ),
        ( "01111001", "10000001", "10100101" ),
        ( "00110011", "10001100", "10100100" ),
        ( "01100001", "11000111", "10110011" ),
        ( "11001011", "01011111", "10111101" ),
        ( "01000010", "00000011", "00111111" ),
        ( "11000001", "10001010", "01110010" ),
        ( "01100110", "00110100", "10110101" ),
        ( "10100010", "00000001", "00100010" ),
        ( "11110001", "00011100", "01000110" ),
        ( "01110101", "11010001", "00111001" ),
        ( "11111101", "01101000", "11101111" ),
        ( "00110101", "01000000", "00111110" ),
        ( "11010111", "10000101", "01111111" ),
        ( "00110011", "00100000", "01101010" ),
        ( "11000111", "10110011", "11011100" ),
        ( "11000111", "01000011", "11001010" ),
        ( "00110011", "00110000", "00000011" ),
        ( "11011100", "01001010", "01000011" ),
        ( "11111100", "10010110", "01101010" ),
        ( "00111011", "01010000", "00100100" ),
        ( "01011110", "11000010", "11010000" ),
        ( "10100100", "00011100", "00000111" ),
        ( "10111111", "11011011", "10101000" ),
        ( "00010001", "11011001", "00100111" ),
        ( "00110110", "01010011", "10010100" ),
        ( "10110101", "10001111", "10000000" ),
        ( "10100110", "11110100", "10110101" ),
        ( "10100000", "11000111", "01001010" ),
        ( "11001010", "01100100", "10111000" ),
        ( "00000101", "00101110", "10110110" ),
        ( "10000100", "10010100", "11101000" ),
        ( "10010101", "00000110", "11110111" ),
        ( "01000111", "00100000", "10101011" ),
        ( "01110100", "11001000", "11110000" ),
        ( "01111010", "10001100", "00111011" ),
        ( "10101011", "01010001", "00101101" ),
        ( "00100010", "11010110", "01110001" ),
        ( "00101001", "01011010", "11101011" ),
        ( "00111100", "11100111", "11111101" ),
        ( "10101100", "00111110", "01011001" ),
        ( "10000110", "10110110", "01101011" ),
        ( "00101101", "00110110", "01011001" ),
        ( "10100111", "01001000", "10110111" ),
        ( "10100111", "10001100", "01110000" ),
        ( "00000000", "11001011", "01100111" ),
        ( "01001000", "01111000", "10011101" ),
        ( "10000011", "10000010", "01011110" ),
        ( "01110011", "10101011", "01010000" ),
        ( "01101000", "00111001", "11101010" ),
        ( "00011011", "10101010", "11000100" ),
        ( "10010101", "01111000", "10111010" ),
        ( "01100011", "10001011", "01011000" ),
        ( "00010010", "10110111", "10111100" ),
        ( "01111110", "10110101", "11000101" ),
        ( "11101000", "00110111", "00010110" ),
        ( "01001010", "10101001", "01000101" ),
        ( "00110101", "01001110", "10110100" ),
        ( "00011100", "00001011", "11111100" ),
        ( "01011100", "01010001", "00101000" ),
        ( "10110001", "01011000", "01001111" ),
        ( "10011011", "01010011", "11000101" ),
        ( "01001100", "00010010", "11100100" ),
        ( "01101111", "01111011", "01000010" ),
        ( "01010111", "01001100", "10000011" ),
        ( "10001001", "10100010", "01001001" ),
        ( "00110001", "11010010", "00010100" ),
        ( "01001001", "01101001", "10111010" ),
        ( "11101001", "01101011", "01100011" ),
        ( "11110001", "00011100", "10001100" ),
        ( "00010100", "11100010", "01111100" ),
        ( "00001110", "11101001", "10010110" ),
        ( "00000010", "11010111", "10111011" ),
        ( "11010101", "01100010", "10011100" ),
        ( "00000000", "10001111", "11100000" ),
        ( "01011111", "00111110", "01111011" ),
        ( "01100101", "00110110", "11000110" ),
        ( "11111110", "11010010", "01001111" ),
        ( "10011110", "01001110", "10010100" ),
        ( "00110001", "10111111", "11010111" ),
        ( "01111001", "01000100", "10000000" ),
        ( "11011110", "11000001", "10010100" ),
        ( "01010011", "01100100", "01111001" ),
        ( "11010010", "10101111", "01001101" ),
        ( "00000100", "10011100", "01001101" ),
        ( "11000001", "11111011", "11111101" ),
        ( "10010111", "11010011", "00110111" ),
        ( "00111000", "01011110", "01100000" ),
        ( "00101011", "11000001", "11001011" ),
        ( "00111010", "01110111", "10001101" ),
        ( "10011000", "10000110", "10111011" ),
        ( "10001011", "01111111", "01100011" ),
        ( "10101001", "01110011", "11110011" ),
        ( "11001101", "01011111", "10111110" ),
        ( "00001111", "11000000", "11110011" ),
        ( "11110101", "11001100", "10100000" ),
        ( "01001111", "00101111", "01110110" ),
        ( "11011000", "00111111", "11010110" ),
        ( "01100001", "11000010", "11001000" ),
        ( "10101001", "11011000", "11000111" ),
        ( "10111100", "00000111", "01010110" ),
        ( "11000111", "10001011", "01101010" ),
        ( "11111001", "10111010", "01011100" ),
        ( "00110010", "00110011", "10011000" ),
        ( "01011100", "10100100", "11000011" ),
        ( "01110111", "01010110", "00110010" ),
        ( "11100011", "11110011", "10000101" ),
        ( "11111100", "11000011", "11010011" ),
        ( "10100110", "10011000", "00110111" ),
        ( "11101010", "01010000", "00001110" ),
        ( "10101100", "00111010", "10001000" ),
        ( "00100111", "01100001", "01100000" ),
        ( "10010001", "11101000", "11010100" ),
        ( "00101100", "00000001", "01011001" ),
        ( "01111010", "10001111", "00011010" ),
        ( "10001011", "10110010", "10111010" ),
        ( "01010110", "11011000", "11111100" ),
        ( "10000100", "01000100", "01101101" ),
        ( "01100110", "00001100", "10010011" ),
        ( "00000110", "01001000", "10100000" ),
        ( "01101100", "11111001", "00110001" ),
        ( "11011110", "00000110", "01110110" ),
        ( "00100001", "00011001", "01110100" ),
        ( "00001101", "11111001", "11111111" ),
        ( "11000001", "01110000", "00101111" ),
        ( "01111000", "00111110", "01111011" ),
        ( "11000110", "11010001", "00011011" ),
        ( "01110001", "01111110", "00011001" ),
        ( "00110101", "10001001", "01001000" ),
        ( "11001011", "00101111", "10101001" ),
        ( "11111100", "10101110", "11000100" ),
        ( "01110001", "01001110", "11111010" ),
        ( "01011011", "01111011", "11111111" ),
        ( "10111100", "11011100", "11100001" ),
        ( "01010000", "01111011", "11000011" ),
        ( "00000000", "10111100", "00011100" ),
        ( "01110011", "01111100", "11100110" ),
        ( "00000011", "11001100", "10000101" ),
        ( "11010001", "01111011", "11111111" ),
        ( "01011000", "01001111", "01011000" ),
        ( "10100001", "00001000", "10111100" ),
        ( "11011011", "11111111", "01111110" ),
        ( "11101011", "11010101", "10110010" ),
        ( "10111110", "01100001", "00001111" ),
        ( "01110011", "01101101", "11000001" ),
        ( "11101010", "00110000", "10010000" ),
        ( "10001000", "01000011", "01011111" ),
        ( "10010111", "11111010", "10011001" ),
        ( "10010010", "10011010", "01011101" ),
        ( "01110010", "01001011", "11100010" ),
        ( "01100100", "11111010", "00010010" ),
        ( "10101011", "11101110", "11101110" ),
        ( "11000110", "00101000", "11110001" ),
        ( "10111000", "00110001", "11001000" ),
        ( "10110000", "11011100", "11011110" ),
        ( "10111000", "00110101", "10010010" ),
        ( "00101111", "10101001", "11111011" ),
        ( "10110100", "10101010", "11010011" ),
        ( "11101011", "11011011", "10010100" ),
        ( "00111010", "10001001", "11000110" ),
        ( "11000001", "00110000", "01110000" ),
        ( "11111011", "10101010", "00011011" ),
        ( "11111100", "10110000", "11000000" ),
        ( "01111000", "01000110", "11101011" ),
        ( "00000000", "00100000", "01010101" ),
        ( "11101001", "11001000", "11001010" ),
        ( "10010010", "10111101", "11101001" ),
        ( "11010010", "01111101", "00111001" ),
        ( "11111101", "00111001", "10011111" ),
        ( "00010001", "11111011", "11101100" ),
        ( "10111111", "00111110", "00001000" ),
        ( "01001001", "01011001", "10100001" ),
        ( "10010000", "11011111", "01001100" ),
        ( "11101001", "10010110", "01110101" ),
        ( "11010011", "10110110", "01001000" ),
        ( "01001110", "10110110", "11111110" ),
        ( "11010111", "10101100", "11000010" ),
        ( "10110001", "10000101", "10010011" ),
        ( "01110110", "10011000", "00000000" ),
        ( "11001111", "11111111", "10000011" ),
        ( "11101110", "00111001", "01100111" ),
        ( "10100011", "11001001", "00110101" ),
        ( "00001001", "00110101", "11101101" ),
        ( "01111111", "01001000", "01100000" ),
        ( "11101111", "00101000", "10000000" ),
        ( "01100001", "00110001", "11011011" ),
        ( "00111101", "11100101", "10110011" ),
        ( "01100101", "10101011", "10110110" ),
        ( "00101100", "01110100", "01001110" ),
        ( "10011010", "01011010", "10011111" ),
        ( "11110011", "01111001", "10010110" ),
        ( "10100111", "11100111", "10111101" ),
        ( "10101011", "11111101", "01100110" ),
        ( "11111110", "11101000", "10000100" ),
        ( "01010110", "11011111", "01110100" ),
        ( "10010111", "00110110", "00110011" ),
        ( "11100010", "01001110", "01010001" ),
        ( "01100101", "00000101", "11111101" ),
        ( "00110111", "00010110", "00000110" ),
        ( "11111110", "01101101", "00000111" ),
        ( "10110011", "10110001", "01100100" ),
        ( "00111010", "00011010", "11000000" ),
        ( "10101000", "01010100", "01010111" ),
        ( "10101000", "01011010", "01000110" ),
        ( "10101010", "01110101", "11100000" ),
        ( "00101100", "11001101", "11001100" ),
        ( "11011011", "01110101", "10000100" ),
        ( "00101111", "01011001", "01000101" ),
        ( "01110101", "01111101", "01001101" ),
        ( "00010111", "00111010", "10111000" ),
        ( "00111100", "10100111", "10110101" ),
        ( "00001011", "00111000", "00001111" ),
        ( "10100011", "00001100", "00010010" ),
        ( "00110000", "01110100", "00111110" ),
        ( "11001100", "01010011", "01011011" ),
        ( "11011010", "01001101", "00010000" ),
        ( "10100001", "11001111", "01011000" ),
        ( "01110000", "00111110", "00000111" ),
        ( "10111111", "01001110", "10101010" ),
        ( "11101100", "11010100", "00000011" ),
        ( "11110001", "00101011", "00100001" ),
        ( "01000010", "00000110", "10110111" ),
        ( "01011001", "01000000", "01011001" ),
        ( "00010010", "10001110", "00011000" ),
        ( "10101011", "11001000", "10100011" ),
        ( "01101111", "00100001", "00111100" ),
        ( "00000101", "01010011", "10011000" ),
        ( "10100110", "10010110", "01101001" ),
        ( "00111001", "01011101", "11101010" ),
        ( "01001000", "01001101", "01010010" ),
        ( "10110110", "00100000", "01010010" ),
        ( "11011101", "10000101", "10011111" ),
        ( "01001110", "10111101", "10101101" ),
        ( "00010101", "01100011", "01011010" ),
        ( "10000010", "11010110", "10100100" ),
        ( "01001100", "11001001", "11100000" ),
        ( "00100111", "00100001", "01110000" ),
        ( "10111101", "01011011", "01011011" ),
        ( "01111100", "10101011", "10011100" ),
        ( "10111001", "01000010", "11111011" ),
        ( "00000101", "10111000", "11011010" ),
        ( "10110111", "10000110", "01011000" ),
        ( "11010001", "10000111", "00110110" ),
        ( "00100011", "00011110", "11010101" ),
        ( "11101010", "01101100", "01010111" ),
        ( "00110000", "00000110", "11010101" ),
        ( "00100101", "11101110", "10010011" ),
        ( "00010100", "11110110", "00010110" ),
        ( "10010010", "11110110", "11110001" ),
        ( "01111101", "10010000", "10100011" ),
        ( "00101111", "00101110", "01111011" ),
        ( "00100101", "00101000", "00001111" ),
        ( "10110100", "00100100", "01101011" ),
        ( "11000010", "01100101", "11110011" ),
        ( "10010011", "11001010", "00010101" ),
        ( "11010001", "01110110", "11101111" ),
        ( "01111010", "01101000", "10011111" ),
        ( "11100011", "10001110", "10011010" ),
        ( "11111111", "00100101", "11100101" ),
        ( "01111101", "11011111", "00100110" ),
        ( "00111101", "10100100", "00011001" ),
        ( "10101011", "01010111", "10100001" ),
        ( "10001000", "01110010", "00000101" ),
        ( "11000111", "10111101", "00011000" ),
        ( "10000101", "00110101", "11110011" ),
        ( "00111010", "00001101", "00010000" ),
        ( "01000101", "11011011", "10100111" ),
        ( "00001111", "00011111", "00000101" ),
        ( "00111111", "00111101", "11110011" ),
        ( "10110011", "11111010", "11111010" ),
        ( "00101101", "11101111", "11001010" ),
        ( "01000011", "01101000", "00111000" ),
        ( "01000000", "00110100", "11100010" ),
        ( "00100110", "10100001", "11001011" ),
        ( "00101101", "01010001", "00111011" ),
        ( "11101111", "00101000", "01101110" ),
        ( "11111001", "10110001", "00101110" ),
        ( "10111011", "00110110", "11010001" ),
        ( "10001101", "10011110", "11001111" ),
        ( "10000100", "00111010", "10001000" ),
        ( "01111100", "01110100", "11000011" ),
        ( "00100000", "01100000", "00001001" ),
        ( "10000100", "10011110", "11011110" ),
        ( "11100111", "00011110", "01110100" ),
        ( "10101111", "10111000", "00100101" ),
        ( "00110100", "00110001", "00101011" ),
        ( "00011001", "10101110", "00000010" ),
        ( "00111100", "10011000", "01011000" ),
        ( "11001110", "10110111", "11010001" ),
        ( "11110100", "01100101", "11110111" ),
        ( "00111100", "01101100", "00010001" ),
        ( "11110100", "10001001", "00000001" ),
        ( "00100110", "01111101", "11010110" ),
        ( "10100100", "11011010", "11000001" ),
        ( "00100100", "10100100", "01010111" ),
        ( "00010100", "00001100", "10001010" ),
        ( "00001111", "11110000", "10101110" ),
        ( "01000010", "01010000", "00111010" ),
        ( "11101011", "01111011", "00011000" ),
        ( "11000111", "11010100", "01001111" ),
        ( "00101010", "00011111", "01100001" ),
        ( "00100111", "01100001", "10000001" ),
        ( "01100111", "11011001", "01000101" ),
        ( "00100111", "11000100", "00010100" ),
        ( "11011100", "11001010", "11011100" ),
        ( "11111110", "11000011", "01101001" ),
        ( "01001010", "00011011", "01111100" ),
        ( "01000111", "11001111", "01110001" ),
        ( "00001010", "00110011", "10001110" ),
        ( "11101010", "10111011", "00001011" ),
        ( "01111100", "11111001", "01000110" ),
        ( "10000011", "00010010", "10000000" ),
        ( "00010101", "00100011", "01000101" ),
        ( "11110010", "11100100", "10001111" ),
        ( "10110111", "10110101", "10001011" ),
        ( "00001011", "00101111", "11001010" ),
        ( "00011000", "00111110", "01000111" ),
        ( "10101111", "00100001", "00110110" ),
        ( "01100100", "10000100", "01011001" ),
        ( "10101101", "11101011", "01101110" ),
        ( "01100000", "10001011", "10110010" ),
        ( "00111001", "11100000", "10101100" ),
        ( "10110101", "01000001", "11010101" ),
        ( "11100010", "00001011", "10010010" ),
        ( "00101100", "00111110", "00011000" ),
        ( "01001110", "10010000", "10001011" ),
        ( "00000011", "01001111", "10000001" ),
        ( "00011100", "01101010", "00001110" ),
        ( "10100110", "11001000", "01010101" ),
        ( "11000011", "01100100", "00110010" ),
        ( "01101001", "11001110", "10101111" ),
        ( "01001110", "01011111", "01010110" ),
        ( "00100000", "00100000", "10110100" ),
        ( "00110000", "01001000", "11000111" ),
        ( "10100001", "00000010", "01000101" ),
        ( "10111011", "01001101", "10101000" ),
        ( "10010010", "01010011", "01000010" ),
        ( "11010110", "00100100", "10001010" ),
        ( "00011101", "11111111", "10110010" ),
        ( "00000010", "10001010", "01110110" )
    );

    constant hsv_data : hsv_array_t := (
        ( "000000000", "11111111", "11111111" ),
        ( "001111000", "11111111", "11111111" ),
        ( "011110000", "11111111", "11111111" ),
        ( "000111100", "11111111", "11111111" ),
        ( "100101100", "11111111", "11111111" ),
        ( "010110100", "11111111", "11111111" ),
        ( "010100001", "10011110", "11110100" ),
        ( "000000011", "11100000", "11110111" ),
        ( "100000110", "00110110", "11100101" ),
        ( "100000101", "10111000", "10011111" ),
        ( "011001000", "11101100", "10010111" ),
        ( "000001000", "01110110", "10100110" ),
        ( "011100011", "11011101", "11101111" ),
        ( "010111010", "10001001", "11110110" ),
        ( "011001000", "11100010", "11111100" ),
        ( "100001110", "10001100", "10000011" ),
        ( "001011100", "10000011", "01101101" ),
        ( "000000000", "10100110", "01110011" ),
        ( "011100100", "00111110", "10100010" ),
        ( "011010011", "11110001", "01110000" ),
        ( "100000001", "01111110", "11011000" ),
        ( "010011100", "00101001", "01111010" ),
        ( "001010000", "11100101", "11011100" ),
        ( "101010111", "01000101", "11100111" ),
        ( "000101101", "11000000", "10110111" ),
        ( "100101000", "10111100", "11000110" ),
        ( "100100100", "11100001", "11111010" ),
        ( "010011110", "11110100", "10100101" ),
        ( "100001011", "10110101", "10010101" ),
        ( "100111111", "11000110", "11000010" ),
        ( "011110101", "11010011", "10000111" ),
        ( "100000100", "01101011", "11110000" ),
        ( "000010011", "01011000", "11110100" ),
        ( "011000011", "10110101", "11010110" ),
        ( "000101000", "10010001", "10100000" ),
        ( "001111010", "10011101", "10000011" ),
        ( "001111000", "01110010", "10100011" ),
        ( "001110100", "10001000", "11001110" ),
        ( "001110100", "11110010", "10101001" ),
        ( "010001011", "11101010", "01100101" ),
        ( "001010100", "11111111", "11100010" ),
        ( "010010101", "11100100", "11000010" ),
        ( "010010101", "11011000", "01010000" ),
        ( "010001010", "11110101", "11010100" ),
        ( "100011100", "11010010", "11000001" ),
        ( "010001111", "11100011", "10111011" ),
        ( "001011000", "11100111", "11101000" ),
        ( "010111100", "11111111", "10101111" ),
        ( "100101111", "11111100", "11110101" ),
        ( "000010011", "00101101", "11110000" ),
        ( "010010100", "00100101", "11110101" ),
        ( "000001110", "10100010", "01111100" ),
        ( "000100100", "10110101", "11100111" ),
        ( "100100100", "10101000", "11100001" ),
        ( "001010000", "01101000", "10111110" ),
        ( "001011010", "01000000", "11110001" ),
        ( "011000011", "10010100", "10011110" ),
        ( "100010111", "11101111", "11100100" ),
        ( "100011111", "10100010", "10010111" ),
        ( "001001001", "11101101", "10010001" ),
        ( "011101100", "01111000", "11000000" ),
        ( "011111011", "10010101", "11100111" ),
        ( "100000000", "10111001", "10011110" ),
        ( "100010011", "11011100", "10110010" ),
        ( "001111000", "01101001", "11001110" ),
        ( "010111010", "10001100", "11110010" ),
        ( "001110000", "11111100", "10101100" ),
        ( "000011111", "10110111", "01001110" ),
        ( "100100101", "10100111", "11111110" ),
        ( "001110101", "10110101", "11011010" ),
        ( "001110100", "01110101", "10111111" ),
        ( "011101011", "11111010", "11111000" ),
        ( "010100001", "10111111", "10101101" ),
        ( "100110000", "01010101", "11010101" ),
        ( "100000010", "10110010", "11011110" ),
        ( "001100001", "11011011", "10111001" ),
        ( "000101111", "11000110", "10011111" ),
        ( "101001000", "10000001", "01000101" ),
        ( "101010001", "11001100", "10101101" ),
        ( "001101000", "11010001", "11110011" ),
        ( "001111000", "00000001", "11101010" ),
        ( "101011010", "01100110", "11010111" ),
        ( "000110001", "01111010", "11001100" ),
        ( "011101111", "10100110", "11110101" ),
        ( "001101001", "10110011", "11001010" ),
        ( "000101111", "11110111", "11001010" ),
        ( "000100001", "10101010", "11001011" ),
        ( "010010101", "01100001", "11110100" ),
        ( "000110101", "01101100", "11001010" ),
        ( "001011001", "11110011", "11111010" ),
        ( "011111010", "11010010", "11101010" ),
        ( "000010101", "11100101", "11111110" ),
        ( "100000100", "11000110", "10111000" ),
        ( "011001010", "11100110", "01101000" ),
        ( "011100001", "11000001", "10111100" ),
        ( "011111100", "01011100", "10001111" ),
        ( "000010100", "11100100", "11101010" ),
        ( "000101110", "10101111", "10010001" ),
        ( "000111011", "10110000", "01110101" ),
        ( "001011011", "11110001", "11110000" ),
        ( "011111100", "10011011", "11101011" ),
        ( "000000010", "11111101", "10001000" ),
        ( "011111011", "01111110", "10011011" ),
        ( "000111110", "11000101", "11001000" ),
        ( "000000000", "10001000", "11100111" ),
        ( "100101111", "10011000", "10110011" ),
        ( "011000000", "00101111", "11100010" ),
        ( "100101110", "11110110", "11110000" ),
        ( "101010001", "10101000", "11101111" ),
        ( "100001100", "10100011", "11101101" ),
        ( "101011100", "00011010", "10001001" ),
        ( "010010111", "10000010", "10111110" ),
        ( "001001110", "10110001", "01111101" ),
        ( "010001010", "10111011", "11101011" ),
        ( "101100100", "10000111", "11100100" ),
        ( "100110010", "01111100", "11101100" ),
        ( "000111000", "10101001", "10101111" ),
        ( "000100110", "11000001", "11110011" ),
        ( "010100001", "11110100", "01100011" ),
        ( "011100010", "11101011", "10000011" ),
        ( "011001011", "00110000", "10101000" ),
        ( "001000101", "11100010", "10110000" ),
        ( "000101100", "10111100", "10101100" ),
        ( "101000010", "11001111", "11111001" ),
        ( "100101011", "11000011", "11110100" ),
        ( "011101011", "11100000", "01101110" ),
        ( "000010001", "00110111", "11000001" ),
        ( "001100011", "11010101", "11001101" ),
        ( "001110000", "01101111", "11001010" ),
        ( "101010010", "11001010", "11000010" ),
        ( "011011001", "11010010", "11100011" ),
        ( "010000100", "11100101", "10110011" ),
        ( "101010011", "00111110", "10111000" ),
        ( "100001011", "01110110", "11111110" ),
        ( "000001001", "10010110", "11011101" ),
        ( "010001010", "11011001", "11100000" ),
        ( "101010001", "01111111", "11110100" ),
        ( "100010000", "00111000", "11011001" ),
        ( "010001011", "10000011", "10101110" ),
        ( "010111100", "11010000", "11010000" ),
        ( "011010010", "01111010", "01111001" ),
        ( "100001101", "01010101", "11010110" ),
        ( "011111001", "11001100", "00111101" ),
        ( "000000000", "01101100", "11001010" ),
        ( "100101110", "11100000", "10011110" ),
        ( "001110100", "10111110", "11001010" ),
        ( "001000100", "10100101", "10011101" ),
        ( "000111110", "11110011", "10011100" ),
        ( "100011010", "11010101", "10111001" ),
        ( "100111010", "00110011", "11100000" ),
        ( "001010010", "01101111", "01010101" ),
        ( "011110001", "11111011", "10001000" ),
        ( "000011101", "10111000", "10110010" ),
        ( "000101100", "00011000", "11101110" ),
        ( "010011001", "11011101", "11110101" ),
        ( "011011010", "00101110", "11101011" ),
        ( "100101001", "01111111", "11101100" ),
        ( "100000001", "11101011", "01010000" ),
        ( "100110011", "11000110", "11111111" ),
        ( "001101010", "11111111", "11100101" ),
        ( "100000100", "00111011", "10000000" ),
        ( "010010111", "11011000", "10100110" ),
        ( "101001010", "10100001", "10101100" ),
        ( "011100101", "01011000", "10100001" ),
        ( "010010000", "01111011", "10111100" ),
        ( "010001100", "00011110", "10011001" ),
        ( "101011100", "10111111", "11100100" ),
        ( "000110110", "11100000", "11110010" ),
        ( "101011110", "10101111", "10001010" ),
        ( "010000001", "10110010", "01100111" ),
        ( "100101001", "10001111", "11000011" ),
        ( "010111111", "10100001", "11100011" ),
        ( "010001111", "01110001", "10000000" ),
        ( "100000110", "11110000", "01001000" ),
        ( "001111011", "10110101", "11101100" ),
        ( "001011000", "00101111", "10001101" ),
        ( "101010111", "11111011", "11001111" ),
        ( "000100001", "01000110", "11110010" ),
        ( "010110100", "10101111", "11101010" ),
        ( "001000110", "01001011", "10111001" ),
        ( "101011001", "11111101", "10101111" ),
        ( "001111001", "11010000", "11100001" ),
        ( "100000010", "01010100", "10111011" ),
        ( "001111011", "10011101", "11111110" ),
        ( "001000101", "11110001", "10010101" ),
        ( "000011010", "10110101", "10011000" ),
        ( "100000011", "11111111", "01011111" ),
        ( "100010110", "10101011", "11011110" ),
        ( "000101011", "11100011", "11110001" ),
        ( "101011100", "10011011", "11001011" ),
        ( "101010100", "11010000", "11011111" ),
        ( "100101101", "11011010", "11000011" ),
        ( "000010111", "11000001", "11101110" ),
        ( "000111011", "11101000", "10101101" ),
        ( "000111000", "11001100", "01111000" ),
        ( "101010010", "11001101", "11011001" ),
        ( "001110101", "11010010", "11000111" ),
        ( "000111000", "11110000", "01111000" ),
        ( "001110001", "10000100", "11000100" ),
        ( "001110001", "11011001", "00110110" ),
        ( "000111001", "11100110", "11100001" ),
        ( "101010010", "10111011", "11011110" ),
        ( "000110111", "11011000", "01110000" ),
        ( "101100011", "11000111", "11001110" ),
        ( "101000000", "00111010", "10111111" ),
        ( "010001001", "10000000", "11101111" ),
        ( "011011010", "11010110", "01101011" ),
        ( "001010101", "10111101", "10000000" ),
        ( "001101011", "11101110", "10100110" ),
        ( "010110001", "01110000", "11000011" ),
        ( "010011111", "01101011", "11101001" ),
        ( "001100001", "01111011", "11000111" ),
        ( "000000111", "11101000", "11001111" ),
        ( "011100100", "01011100", "10100000" ),
        ( "001010011", "01011000", "11110010" ),
        ( "101001010", "01100101", "11110100" ),
        ( "001110000", "10011111", "01100011" ),
        ( "011100011", "00111101", "11101011" ),
        ( "011100011", "11010100", "10111111" ),
        ( "010111011", "11101010", "10100010" ),
        ( "011100000", "00101111", "11110011" ),
        ( "000001010", "11101110", "10110101" ),
        ( "011010110", "10010010", "11001110" ),
        ( "000111111", "11111101", "11101001" ),
        ( "011000100", "10011011", "10010101" ),
        ( "001011010", "11000001", "11110001" ),
        ( "011001010", "11111001", "11111110" ),
        ( "001101001", "00100010", "11001110" ),
        ( "100011101", "01101111", "11101010" ),
        ( "011100100", "11001010", "11000100" ),
        ( "000001111", "11010011", "01101001" ),
        ( "011100100", "10010001", "10110110" ),
        ( "001111000", "11000110", "11011100" ),
        ( "010100000", "11100011", "11011101" ),
        ( "101011111", "01101010", "11011111" ),
        ( "100101001", "00011001", "11110010" ),
        ( "011101011", "10011001", "11101110" ),
        ( "001011010", "10110111", "10000111" ),
        ( "001101010", "10110101", "11111010" ),
        ( "001110001", "11100001", "11000110" ),
        ( "100101011", "10101000", "11110111" ),
        ( "000000111", "10110100", "11001010" ),
        ( "000001110", "11111000", "11000001" ),
        ( "011000011", "01011001", "11010000" ),
        ( "100001110", "01111100", "11011011" ),
        ( "010100011", "10110001", "10011110" ),
        ( "010100001", "11110001", "11001100" ),
        ( "000000110", "10110010", "10010110" ),
        ( "101010000", "11001010", "11110000" ),
        ( "011000000", "10100100", "11101011" ),
        ( "100001011", "10100001", "11101110" ),
        ( "001111110", "10010100", "10100011" ),
        ( "011001100", "11011101", "11110010" ),
        ( "010001111", "01110001", "11001101" ),
        ( "011100010", "10000110", "11010001" ),
        ( "001110100", "10010001", "11000110" ),
        ( "001111101", "00111010", "10110011" ),
        ( "100111100", "11001101", "11101101" ),
        ( "000000100", "10000011", "11001010" ),
        ( "011111111", "01011000", "10000101" ),
        ( "010001111", "11110100", "11001010" ),
        ( "001100011", "10101101", "01011000" ),
        ( "000011011", "11000011", "11010111" ),
        ( "010011101", "01100001", "11011110" ),
        ( "000000100", "00111010", "10110010" ),
        ( "101001100", "11111000", "11100110" ),
        ( "100110100", "10010110", "10000110" ),
        ( "001111011", "11101000", "11001100" ),
        ( "001000010", "01100101", "11101000" ),
        ( "100111100", "11110011", "01010111" ),
        ( "011111010", "01110010", "10100000" ),
        ( "011100010", "00011111", "11101101" ),
        ( "011101101", "10100001", "11111010" ),
        ( "011101101", "11011101", "11111010" ),
        ( "011111000", "10010010", "11011100" ),
        ( "101000010", "01100010", "11110110" ),
        ( "000101011", "11111010", "11101100" ),
        ( "001111011", "11001110", "10011101" ),
        ( "011111110", "10001001", "01001100" ),
        ( "010001110", "10101100", "01100110" ),
        ( "000010010", "11110000", "11111111" ),
        ( "000010111", "11110100", "10010100" ),
        ( "001111111", "11110001", "11010011" ),
        ( "100000101", "10001010", "11111110" ),
        ( "001100011", "01110001", "11111101" ),
        ( "000010110", "01101001", "10011001" ),
        ( "101100001", "11101111", "11110111" ),
        ( "011100100", "10100110", "01010100" ),
        ( "001111011", "11010001", "01110110" ),
        ( "101001100", "11011011", "11001001" ),
        ( "011001111", "01111001", "01111010" ),
        ( "001101010", "11111111", "10111110" ),
        ( "011111101", "01111001", "11011001" ),
        ( "010001101", "11001011", "11010101" ),
        ( "001011001", "01110111", "11011110" ),
        ( "100100000", "11010110", "10111000" ),
        ( "000010100", "11100101", "10011101" ),
        ( "011101001", "10000101", "11001000" ),
        ( "000000110", "11110010", "11011011" ),
        ( "010100000", "01110001", "11111001" ),
        ( "000110100", "11111100", "11111000" ),
        ( "010010000", "11101011", "10011110" ),
        ( "000010100", "11001101", "11011010" ),
        ( "011011010", "01111111", "00111100" ),
        ( "000001111", "11101011", "10011010" ),
        ( "100010011", "11100100", "11010110" ),
        ( "011110011", "11111001", "10000100" ),
        ( "011100000", "10100011", "10001100" ),
        ( "001011100", "11111010", "10110111" ),
        ( "100001110", "01001001", "11101011" ),
        ( "100000001", "11100000", "10000111" ),
        ( "010100010", "01000110", "10010100" ),
        ( "100010110", "11000011", "11001100" ),
        ( "001010001", "11101000", "11001000" ),
        ( "101001011", "10100110", "11100100" ),
        ( "010010111", "01110010", "11111011" ),
        ( "001111000", "10101101", "10111100" ),
        ( "100110011", "10010101", "11000010" ),
        ( "011001101", "11101000", "10010011" ),
        ( "101100000", "01101110", "11110001" ),
        ( "011010110", "10011100", "00110001" ),
        ( "001100100", "10100011", "01110010" ),
        ( "101001010", "11011110", "11011110" ),
        ( "001101000", "11000100", "11111011" ),
        ( "011011101", "11110010", "11110000" ),
        ( "010110111", "01010001", "11111101" ),
        ( "101001111", "10010100", "11100001" ),
        ( "001101001", "10011001", "10011001" ),
        ( "011100000", "11001010", "11000001" ),
        ( "001100001", "01011111", "11001001" ),
        ( "010000110", "10011000", "11010101" ),
        ( "000010010", "10110101", "10110001" ),
        ( "100000111", "11011010", "11001001" ),
        ( "010110100", "11100011", "10001101" ),
        ( "101000000", "10110111", "11001110" ),
        ( "101001000", "11000100", "11101110" ),
        ( "101100010", "11101110", "11100110" ),
        ( "010101000", "11011110", "11000101" ),
        ( "010000110", "11110001", "10111100" ),
        ( "001001111", "11101101", "11001110" ),
        ( "000010000", "01111101", "10100000" ),
        ( "001001010", "11010110", "11110101" ),
        ( "011001001", "11101001", "11111010" ),
        ( "011111010", "10100111", "10101011" ),
        ( "100111100", "11101011", "11100100" ),
        ( "011111101", "11010110", "11101000" ),
        ( "101000111", "01011111", "10100000" ),
        ( "011111001", "10111010", "10111111" ),
        ( "001111011", "01011101", "10110111" ),
        ( "011100100", "01110111", "11111100" ),
        ( "100001011", "01011000", "11000001" ),
        ( "100101000", "01111000", "10111000" ),
        ( "100100110", "11110011", "11001100" ),
        ( "010100001", "10000010", "11101000" ),
        ( "011100110", "11010011", "10101010" ),
        ( "101000111", "11110101", "10000100" ),
        ( "000111010", "11000000", "01001001" ),
        ( "001110001", "11001001", "11111110" ),
        ( "101000110", "11000111", "01101110" ),
        ( "011001000", "01011010", "11100100" ),
        ( "100101000", "11010011", "10010100" ),
        ( "001001111", "01111110", "11010011" ),
        ( "010110101", "10001000", "11110001" ),
        ( "000111111", "10101000", "11100110" ),
        ( "000010111", "10010011", "11010001" ),
        ( "101010000", "11110100", "11111001" ),
        ( "010100000", "11000100", "11101110" ),
        ( "011000111", "11011001", "10100010" ),
        ( "000011000", "01111001", "01111010" ),
        ( "000111110", "10111011", "11110000" ),
        ( "101100110", "11011101", "11100111" ),
        ( "100101000", "11000001", "01110100" ),
        ( "001011000", "01010010", "10010101" ),
        ( "001000001", "10111011", "10111101" ),
        ( "101001111", "11110010", "11001011" ),
        ( "001010000", "10110110", "11010010" ),
        ( "011011110", "11000001", "10101111" ),
        ( "011101010", "11111100", "01100000" ),
        ( "000110110", "11010010", "10110110" ),
        ( "000010000", "11110110", "00111100" ),
        ( "010101111", "11101110", "11000110" ),
        ( "010010011", "00101100", "10010110" ),
        ( "000100100", "01001111", "10011110" ),
        ( "100001110", "01111101", "01001101" ),
        ( "011010111", "10101110", "11100010" ),
        ( "000010101", "11001011", "01101101" ),
        ( "000010010", "10010010", "01110101" ),
        ( "001000101", "10100011", "11010100" ),
        ( "100111111", "11010111", "11111000" ),
        ( "101000111", "11011001", "10101000" ),
        ( "100101100", "10000110", "01001010" ),
        ( "011111111", "01110010", "01000101" ),
        ( "010011000", "11111100", "11101100" ),
        ( "101011001", "10100011", "10111110" ),
        ( "100100011", "11111000", "10111000" ),
        ( "001011001", "10010100", "10010101" ),
        ( "010000001", "11111101", "11110001" ),
        ( "000011000", "01100001", "01100001" ),
        ( "010000001", "11100111", "10011001" ),
        ( "011110111", "10010100", "11101010" ),
        ( "000010010", "01101001", "10001100" ),
        ( "011010000", "11010000", "01111111" ),
        ( "010100010", "11011111", "11000011" ),
        ( "011101101", "11010111", "11010110" ),
        ( "100100111", "11011101", "10110111" ),
        ( "011011100", "10100111", "01100011" ),
        ( "011110111", "01010000", "01101000" ),
        ( "010110101", "10111010", "11010011" ),
        ( "100010111", "10011010", "11000101" ),
        ( "101011010", "10110010", "10101110" ),
        ( "001111111", "00100000", "10110110" ),
        ( "101001000", "00111000", "10111001" ),
        ( "000111010", "01100110", "11000011" ),
        ( "011010110", "10101000", "10110001" ),
        ( "010010100", "11110001", "10011011" ),
        ( "011110100", "10100101", "11101110" ),
        ( "001000000", "10001110", "11110111" ),
        ( "011111111", "11101011", "11110111" ),
        ( "001110011", "10100111", "11100110" ),
        ( "000010010", "01010101", "01111110" ),
        ( "000110110", "10010110", "11010010" ),
        ( "011011110", "10100110", "11101110" ),
        ( "001011111", "01111001", "10010111" ),
        ( "100101110", "11010111", "11111101" ),
        ( "101000110", "11001111", "11000000" ),
        ( "000111011", "10101110", "11010100" ),
        ( "001011000", "11111010", "10101111" ),
        ( "000011100", "11010110", "10101111" ),
        ( "100101001", "10110101", "10110000" ),
        ( "000010110", "10011110", "11011111" ),
        ( "011101011", "10001100", "10100101" ),
        ( "000011101", "11110011", "11011001" ),
        ( "001110100", "01101000", "10001011" ),
        ( "000101111", "10101100", "10110100" ),
        ( "011011111", "11100000", "10101110" ),
        ( "010001010", "11111111", "11110100" ),
        ( "000010001", "00100011", "11100000" ),
        ( "000110110", "11100011", "10101110" ),
        ( "011111111", "01101101", "11010100" ),
        ( "000101011", "11110101", "11110011" ),
        ( "011111011", "10011101", "11101001" ),
        ( "100001100", "01101010", "10010100" ),
        ( "101011110", "11010100", "11010010" ),
        ( "010111111", "11011110", "11000011" ),
        ( "001011111", "10110001", "10000000" ),
        ( "011101111", "10001001", "11001111" ),
        ( "000110111", "11011001", "11010100" ),
        ( "000001101", "11001011", "11111011" ),
        ( "000100001", "10010011", "11101000" ),
        ( "011001011", "01010010", "01000001" ),
        ( "001101101", "10101011", "10101011" ),
        ( "010100011", "11011111", "10100100" ),
        ( "001101001", "10011000", "11111111" ),
        ( "000011001", "11011100", "11100110" ),
        ( "000100110", "11101100", "11010001" ),
        ( "101000111", "10101101", "11010111" ),
        ( "011100110", "11111111", "10000101" ),
        ( "011100101", "11101111", "11100000" ),
        ( "001101011", "11101101", "10000101" ),
        ( "011100010", "11111110", "11111111" ),
        ( "100111100", "10111000", "10000010" ),
        ( "001111000", "11110010", "11111101" ),
        ( "100100111", "11000110", "11110001" ),
        ( "011110100", "11011000", "10011010" ),
        ( "011010010", "11000010", "00111011" ),
        ( "000011010", "10101010", "11011010" ),
        ( "100000000", "10110110", "10110100" ),
        ( "011101100", "10010010", "11101011" ),
        ( "100011000", "01111010", "11111000" ),
        ( "101000110", "11010100", "11101110" ),
        ( "001010101", "10000110", "10111000" ),
        ( "001100000", "10000000", "11101100" ),
        ( "000110011", "11101011", "11101010" ),
        ( "000011000", "11111010", "01100111" ),
        ( "000100001", "10110011", "11001000" ),
        ( "101010010", "10010010", "10110011" ),
        ( "001101101", "10101110", "11011010" ),
        ( "001010100", "10100100", "10100100" ),
        ( "101001001", "11011010", "11111010" ),
        ( "000010001", "00110101", "11100100" ),
        ( "100010011", "11111111", "10111011" ),
        ( "011011010", "11010110", "11001010" ),
        ( "000000010", "11001010", "10111111" ),
        ( "100101101", "01010010", "11011011" ),
        ( "000100001", "10001111", "11100011" ),
        ( "101011011", "11011011", "11111001" ),
        ( "101001011", "10111100", "01101100" ),
        ( "010001100", "01100100", "11110111" ),
        ( "101001010", "11011100", "11111001" ),
        ( "000001100", "11011010", "10000011" ),
        ( "000010001", "11111010", "01101001" ),
        ( "100011000", "11010101", "11111111" ),
        ( "011001001", "10101010", "11001011" ),
        ( "010100000", "01101100", "11011101" ),
        ( "100110110", "10010111", "11010100" ),
        ( "001111101", "11010101", "11010001" ),
        ( "000100010", "11111011", "11101110" ),
        ( "001100001", "01100010", "11010100" ),
        ( "011111101", "11001000", "11011010" ),
        ( "100000001", "01001001", "11001110" ),
        ( "011111010", "11100100", "11010111" ),
        ( "101000011", "11100101", "01111010" ),
        ( "100000000", "11010011", "10101011" ),
        ( "010011111", "11010111", "11110110" ),
        ( "100100111", "11110101", "00111000" ),
        ( "101100001", "01011001", "10100011" ),
        ( "101000111", "01111100", "11111000" ),
        ( "100111010", "01110101", "11100001" ),
        ( "000110010", "10011101", "10111100" ),
        ( "010010010", "10011101", "01110000" ),
        ( "001110100", "01111101", "11001110" ),
        ( "000111011", "11110100", "11110011" ),
        ( "101010100", "10010101", "10110110" ),
        ( "011110101", "01101110", "01101100" ),
        ( "100001010", "11100110", "01010011" ),
        ( "011110000", "10110000", "10001000" ),
        ( "011011010", "01001001", "11000010" ),
        ( "010111100", "11010110", "11100001" ),
        ( "011011011", "10101011", "10100100" ),
        ( "011000100", "11101110", "11110010" ),
        ( "000000101", "01011100", "11100010" ),
        ( "011100011", "10010100", "10110100" ),
        ( "101100010", "11011011", "10100100" ),
        ( "100100101", "10001011", "00110101" ),
        ( "000011100", "10000111", "10100100" ),
        ( "100110100", "10000101", "11010000" ),
        ( "010110001", "11101010", "11001111" ),
        ( "101001000", "11100000", "10110101" ),
        ( "011111011", "11100100", "10100010" ),
        ( "011101010", "11010010", "11000001" ),
        ( "001100000", "10010000", "11001101" ),
        ( "001101110", "11011001", "01011001" ),
        ( "100101000", "10001010", "11010100" ),
        ( "101100011", "01101111", "11101011" ),
        ( "001011010", "01001100", "10111111" ),
        ( "100011110", "00011100", "01010001" ),
        ( "101100011", "01101100", "10001011" ),
        ( "010101100", "10110001", "11001011" ),
        ( "000101001", "11101011", "11011011" ),
        ( "100110011", "11011000", "11111001" ),
        ( "010101010", "11100111", "11000011" ),
        ( "010001011", "11111010", "11111101" ),
        ( "010000011", "11000100", "11011011" ),
        ( "011010001", "11111111", "11001100" ),
        ( "000110010", "10000011", "11111001" ),
        ( "011111110", "01110001", "11111101" ),
        ( "010111101", "11111010", "11110100" ),
        ( "011110000", "01101010", "10011110" ),
        ( "011001010", "11000010", "11111011" ),
        ( "010000100", "11111111", "10100000" ),
        ( "011011101", "11010011", "11101000" ),
        ( "010101100", "11100000", "11111010" ),
        ( "000101001", "01110101", "11110101" ),
        ( "010110111", "00101111", "10011011" ),
        ( "100001010", "11111010", "10101101" ),
        ( "100110000", "11111100", "11000001" ),
        ( "010000101", "01010000", "10001000" ),
        ( "001011100", "01110000", "11000101" ),
        ( "011000100", "00111101", "11000010" ),
        ( "100010111", "10010011", "11011101" ),
        ( "010110000", "11100100", "00010011" ),
        ( "011111010", "10010001", "11011010" ),
        ( "001111001", "01011100", "10100101" ),
        ( "010110111", "11011001", "10111111" ),
        ( "100000110", "01110001", "01100111" ),
        ( "000100110", "00110111", "11011000" ),
        ( "001101111", "00011100", "10110110" ),
        ( "100110000", "10100001", "11111000" ),
        ( "100000010", "11011001", "01011110" ),
        ( "100001001", "11110110", "10110100" ),
        ( "000001100", "10010111", "11101001" ),
        ( "011110100", "10100110", "11010101" ),
        ( "011110111", "11111111", "11011011" ),
        ( "100010010", "01000111", "10110110" ),
        ( "001011101", "11100010", "01100100" ),
        ( "000001001", "01011010", "11100011" ),
        ( "100001010", "11010000", "11001101" ),
        ( "100111001", "11111010", "01101011" ),
        ( "101011100", "11010111", "11000111" ),
        ( "101100100", "11001101", "11000101" ),
        ( "001010010", "01010001", "11000110" ),
        ( "010001111", "11010101", "11011110" ),
        ( "011100111", "10110101", "11001001" ),
        ( "000010000", "11011010", "10011000" ),
        ( "100110011", "10010110", "01101001" ),
        ( "011000011", "10101010", "10100000" ),
        ( "100110101", "01110001", "11011101" ),
        ( "001011100", "01001000", "11011111" ),
        ( "010101001", "11000101", "10101000" ),
        ( "000011001", "11000010", "01101110" ),
        ( "100011011", "10100010", "01100110" ),
        ( "000000000", "11011110", "11110000" ),
        ( "001010101", "10101111", "11101000" ),
        ( "100101111", "11101100", "10110000" ),
        ( "000010010", "01100010", "01101101" ),
        ( "011001000", "11111011", "11111100" ),
        ( "001001000", "11101011", "01111000" ),
        ( "100100011", "11110010", "11111011" ),
        ( "011111111", "11011000", "10110101" ),
        ( "000100100", "11011001", "11111001" ),
        ( "010000001", "10010000", "10010110" ),
        ( "000110010", "11000010", "11110001" ),
        ( "011011011", "01010011", "11100011" ),
        ( "010100101", "10101010", "11011110" ),
        ( "101010001", "10011001", "10010010" ),
        ( "100011000", "10110011", "11000100" ),
        ( "001001101", "01101010", "01111111" ),
        ( "100001010", "11110010", "11110101" ),
        ( "010110001", "00110010", "01100101" ),
        ( "000000110", "10000110", "10100101" ),
        ( "000001011", "01111111", "11101010" ),
        ( "000010011", "10000001", "10111111" ),
        ( "011100101", "01001001", "11011101" ),
        ( "001110100", "11010111", "10111010" ),
        ( "011111101", "11001001", "11111101" ),
        ( "001101101", "11001011", "11101111" ),
        ( "001100001", "11011101", "11111000" ),
        ( "010000100", "01100110", "11100010" ),
        ( "100101111", "11100010", "11001100" ),
        ( "001001010", "11110111", "10100111" ),
        ( "000111000", "10011101", "10110111" ),
        ( "101100001", "11111100", "11101010" ),
        ( "100000110", "10000101", "01101101" ),
        ( "010101111", "10101000", "11010100" ),
        ( "001110001", "10111001", "11100111" ),
        ( "000111111", "11111100", "11111001" ),
        ( "010000011", "11011011", "01100101" ),
        ( "011110000", "11010110", "11011100" ),
        ( "001000111", "11001010", "11110100" ),
        ( "011101100", "01100011", "11011101" ),
        ( "100101010", "11110100", "01111001" ),
        ( "010100111", "10111110", "10100010" ),
        ( "010000111", "11000001", "00111110" ),
        ( "001110001", "11011101", "11101010" ),
        ( "010110010", "10001010", "11011010" ),
        ( "010100001", "11000011", "11011001" ),
        ( "011100010", "10111001", "10100001" ),
        ( "100000000", "10010011", "11010111" ),
        ( "100110110", "10101110", "11011110" ),
        ( "100101010", "10111001", "10001100" ),
        ( "001001000", "11000111", "11111011" ),
        ( "100000010", "10100001", "10111110" ),
        ( "101010000", "00111100", "11100110" ),
        ( "000010010", "10100101", "10100011" ),
        ( "101001100", "10110111", "10111101" ),
        ( "101001110", "01010111", "10100110" ),
        ( "101011110", "10111000", "10011011" ),
        ( "011001001", "11000001", "11000011" ),
        ( "011001100", "10001011", "10111010" ),
        ( "000000001", "01001101", "10001101" ),
        ( "100001000", "01101110", "11000100" ),
        ( "000110001", "11111111", "01100110" ),
        ( "100010100", "10000100", "11111011" ),
        ( "100010110", "10100100", "11010110" ),
        ( "010000101", "10001111", "11111010" ),
        ( "001101010", "10000110", "11110011" ),
        ( "011100001", "10111100", "11101100" ),
        ( "010101001", "10101111", "11011000" ),
        ( "000011110", "10111101", "11000011" ),
        ( "101001101", "11011011", "11011111" ),
        ( "010000001", "01100100", "10000110" ),
        ( "011100110", "01000100", "10100101" ),
        ( "011000001", "10101111", "10100100" ),
        ( "010101000", "10000010", "11000111" ),
        ( "100110100", "10000111", "11001011" ),
        ( "100101111", "11110011", "01000010" ),
        ( "000010010", "01101000", "11000001" ),
        ( "100000111", "10110101", "10110101" ),
        ( "101011100", "11111101", "10100010" ),
        ( "101011101", "11100001", "11110001" ),
        ( "001100001", "10111001", "11010001" ),
        ( "100110010", "10010110", "11111101" ),
        ( "010101001", "00101011", "01000000" ),
        ( "000000100", "01101000", "11010111" ),
        ( "011111111", "10110010", "01101010" ),
        ( "100001101", "00101111", "11011100" ),
        ( "100101010", "10101010", "11001010" ),
        ( "000111000", "11110000", "00110011" ),
        ( "000000010", "10110001", "11011100" ),
        ( "000010010", "10010011", "11111100" ),
        ( "001011001", "10001100", "01010000" ),
        ( "010111100", "10001011", "11010000" ),
        ( "000001000", "11110100", "10100100" ),
        ( "001011101", "00111011", "11011011" ),
        ( "001111110", "11101011", "11011001" ),
        ( "011011110", "10100001", "10010100" ),
        ( "000010000", "01001010", "10110101" ),
        ( "010000011", "01010001", "11110100" ),
        ( "001001111", "10100000", "11000111" ),
        ( "100110111", "10000000", "11001010" ),
        ( "011100011", "11110111", "10110110" ),
        ( "011100111", "01101101", "11101000" ),
        ( "100010011", "11111000", "11110111" ),
        ( "100000000", "11001111", "10101011" ),
        ( "011001000", "10000011", "11110000" ),
        ( "001001010", "10010011", "10001100" ),
        ( "000010001", "10111011", "10101011" ),
        ( "010010010", "11010110", "11010110" ),
        ( "011100001", "11010010", "11101011" ),
        ( "010111011", "11000010", "11111101" ),
        ( "101011010", "10100011", "10101100" ),
        ( "001100011", "01101001", "10110110" ),
        ( "011100100", "01111110", "01011001" ),
        ( "100100011", "10011010", "10110111" ),
        ( "000011110", "01010011", "10100111" ),
        ( "010010110", "11111111", "11001011" ),
        ( "011001111", "10001010", "10011101" ),
        ( "000111010", "01001000", "10000011" ),
        ( "001100001", "10000111", "10101011" ),
        ( "011111111", "11000000", "11101010" ),
        ( "010111110", "11011011", "11000100" ),
        ( "100001010", "01011010", "10111010" ),
        ( "001101100", "01011101", "10001011" ),
        ( "010110110", "11100110", "10111100" ),
        ( "011000010", "01011011", "11000101" ),
        ( "000001001", "11100110", "11101000" ),
        ( "001110101", "10010110", "10101001" ),
        ( "011100101", "10110011", "10110100" ),
        ( "011110100", "11110011", "11111100" ),
        ( "000101111", "10010000", "01011100" ),
        ( "000000101", "10001101", "10110001" ),
        ( "100010101", "10010011", "11000101" ),
        ( "100000000", "11101010", "11100100" ),
        ( "001001001", "01110110", "01111011" ),
        ( "011111100", "01101011", "10000011" ),
        ( "001001101", "10001100", "10100010" ),
        ( "001101111", "11100110", "11010010" ),
        ( "011100000", "10011010", "10111010" ),
        ( "000000011", "10010010", "11101001" ),
        ( "101001001", "11100001", "11110001" ),
        ( "010010110", "11101000", "11100010" ),
        ( "010011101", "11101111", "11101001" ),
        ( "010101100", "11111100", "11010111" ),
        ( "101001010", "10001001", "11010101" ),
        ( "011001010", "11111111", "11100000" ),
        ( "100010000", "01111110", "01111011" ),
        ( "100000011", "10111001", "11000110" ),
        ( "000101100", "10101111", "11111110" ),
        ( "100110100", "10000001", "10011110" ),
        ( "010111101", "11000100", "11010111" ),
        ( "100100101", "01110111", "10000000" ),
        ( "000100100", "01010101", "11011110" ),
        ( "011010110", "01010000", "01111001" ),
        ( "000101100", "10100001", "11010010" ),
        ( "010010100", "11111000", "10011100" ),
        ( "010110110", "00111100", "11111101" ),
        ( "001010100", "10111100", "11010011" ),
        ( "010110111", "01101010", "01100000" ),
        ( "010111000", "11001000", "11001011" ),
        ( "011000100", "10010110", "10001101" ),
        ( "100000100", "01001000", "10111011" ),
        ( "000101010", "01001001", "10001011" ),
        ( "100001001", "10000110", "11110011" ),
        ( "100110101", "10001000", "11001101" ),
        ( "011000010", "11101111", "11110011" ),
        ( "000011111", "01011000", "11110101" ),
        ( "100001011", "10011001", "01110110" ),
        ( "100101101", "10110100", "11011000" ),
        ( "010111000", "10000011", "11001000" ),
        ( "010011110", "00110111", "11011000" ),
        ( "101001110", "11110101", "10111100" ),
        ( "000010101", "01110111", "11000111" ),
        ( "000100011", "10100000", "11111001" ),
        ( "011110000", "10101011", "10011000" ),
        ( "011000111", "10000110", "11000011" ),
        ( "000011111", "10010011", "01110111" ),
        ( "001000101", "01110011", "11110011" ),
        ( "101011000", "00111001", "11111100" ),
        ( "000110100", "10101010", "10100110" ),
        ( "000010010", "11101111", "11101010" ),
        ( "100111111", "10101001", "10101100" ),
        ( "010110010", "10011000", "01100001" ),
        ( "010100110", "01011111", "11101000" ),
        ( "100001101", "11111100", "01011001" ),
        ( "001000111", "11010000", "10001111" ),
        ( "010111111", "01000000", "10111010" ),
        ( "011000010", "10100111", "11111100" ),
        ( "101000010", "01111011", "10000100" ),
        ( "100011000", "11101010", "10010011" ),
        ( "011010111", "11110101", "10100000" ),
        ( "001100111", "11001100", "11111001" ),
        ( "101001001", "11111000", "11011110" ),
        ( "011110101", "11001000", "01110100" ),
        ( "010110110", "11110010", "11111111" ),
        ( "000011010", "11000000", "11000001" ),
        ( "100101001", "01111110", "01111011" ),
        ( "001000000", "11011110", "11010001" ),
        ( "001000100", "11001100", "01111110" ),
        ( "010000101", "10011100", "10001001" ),
        ( "100111010", "11000011", "11001011" ),
        ( "101011000", "01001110", "11111100" ),
        ( "011111100", "10101111", "11111010" ),
        ( "011100101", "10100100", "11111111" ),
        ( "010111101", "00101001", "11100001" ),
        ( "011011010", "10010110", "11000011" ),
        ( "010000000", "11111111", "10111100" ),
        ( "011101100", "01111111", "11100110" ),
        ( "010011110", "11111011", "11001100" ),
        ( "100010111", "10000100", "11111111" ),
        ( "100101100", "00011010", "01011000" ),
        ( "100100011", "11110100", "10111100" ),
        ( "001001101", "10000001", "11111111" ),
        ( "000100100", "00111101", "11101011" ),
        ( "000011100", "11101010", "10111110" ),
        ( "011110100", "01101110", "11000001" ),
        ( "101001010", "11001010", "11101010" ),
        ( "101010000", "10000001", "10001000" ),
        ( "001111001", "01100100", "11111010" ),
        ( "001000100", "01100101", "10011010" ),
        ( "011111111", "10101010", "11100010" ),
        ( "001100011", "11101100", "11111010" ),
        ( "010110100", "01000111", "11101110" ),
        ( "100011111", "11010100", "11110001" ),
        ( "100100101", "11000000", "11001000" ),
        ( "010110111", "00110100", "11011110" ),
        ( "100111110", "10110101", "10111000" ),
        ( "011001101", "11001111", "11111011" ),
        ( "011111110", "00110001", "11010011" ),
        ( "000110000", "01011110", "11101011" ),
        ( "011001111", "10110100", "11000110" ),
        ( "101001110", "10111111", "11000001" ),
        ( "000100110", "11100011", "11111011" ),
        ( "101011100", "01001100", "11111100" ),
        ( "100000010", "10110011", "11101011" ),
        ( "011011010", "11111111", "01010101" ),
        ( "101100101", "00100100", "11101001" ),
        ( "011010011", "01011111", "11101001" ),
        ( "000011010", "10111001", "11010010" ),
        ( "101001001", "11000101", "11111101" ),
        ( "010110000", "11101101", "11111011" ),
        ( "000010001", "11110100", "10111111" ),
        ( "011100110", "10001011", "10100001" ),
        ( "001011101", "10101000", "11011111" ),
        ( "000010001", "01111110", "11101001" ),
        ( "000101111", "10100111", "11010011" ),
        ( "011001101", "10110000", "11111110" ),
        ( "101001010", "00110011", "11010111" ),
        ( "101010101", "00111111", "10110001" ),
        ( "001001010", "11111111", "10011000" ),
        ( "001010100", "01111100", "11111111" ),
        ( "101011001", "11000001", "11101110" ),
        ( "001001100", "10111011", "11001001" ),
        ( "011100101", "11110101", "11101101" ),
        ( "101001110", "01101110", "01111111" ),
        ( "101001110", "11010100", "11101111" ),
        ( "100000000", "11000101", "11011011" ),
        ( "010100010", "10111011", "11100101" ),
        ( "010111101", "01110001", "10110110" ),
        ( "010010100", "10011110", "01110100" ),
        ( "100100111", "01101110", "10011111" ),
        ( "101011010", "10000000", "11110011" ),
        ( "010001100", "01000110", "11100111" ),
        ( "001011101", "10011000", "11111101" ),
        ( "000110001", "01111010", "11111110" ),
        ( "010000101", "10011100", "11011111" ),
        ( "000000001", "10101000", "10010111" ),
        ( "101100111", "10100110", "11100010" ),
        ( "100000111", "11111001", "11111101" ),
        ( "000010011", "11100011", "00110111" ),
        ( "000011000", "11110111", "11111110" ),
        ( "000111010", "01110000", "10110011" ),
        ( "011111011", "11011100", "11000000" ),
        ( "101100110", "01111111", "10101000" ),
        ( "000001100", "10010100", "10101000" ),
        ( "100001101", "01111001", "11100000" ),
        ( "010110011", "11001000", "11001101" ),
        ( "101100000", "01110110", "11011011" ),
        ( "010010111", "01111000", "01011001" ),
        ( "001000110", "01100001", "01111101" ),
        ( "011100011", "11011111", "10111000" ),
        ( "010111011", "10101010", "10110101" ),
        ( "001111101", "11001100", "00111000" ),
        ( "101100110", "11101100", "10100011" ),
        ( "010000100", "10010101", "01110100" ),
        ( "101100101", "10010111", "11001100" ),
        ( "000010010", "11101100", "11011010" ),
        ( "001010100", "10010010", "11001111" ),
        ( "000011111", "11101111", "01110000" ),
        ( "100111000", "10010110", "10111111" ),
        ( "000110101", "11111011", "11101100" ),
        ( "000000010", "11011100", "11110001" ),
        ( "100000100", "11110110", "10110111" ),
        ( "100101100", "01000111", "01011001" ),
        ( "001111010", "11011110", "10001110" ),
        ( "001101100", "00101111", "11001000" ),
        ( "101010100", "10110011", "01101111" ),
        ( "011010001", "11110110", "10011000" ),
        ( "000101100", "01011101", "10100110" ),
        ( "011100100", "11000000", "11101010" ),
        ( "011010010", "00011111", "01010010" ),
        ( "101010100", "11010010", "10110110" ),
        ( "101010111", "01100101", "11011101" ),
        ( "010101011", "10010101", "10111101" ),
        ( "010101101", "11001000", "01100011" ),
        ( "010010000", "01100100", "11010110" ),
        ( "010111110", "10101000", "11100000" ),
        ( "011110100", "10110011", "01110000" ),
        ( "000000000", "10000100", "10111101" ),
        ( "010100000", "01000110", "10101011" ),
        ( "100010110", "10111011", "11111011" ),
        ( "010111110", "11111001", "11011010" ),
        ( "000011101", "10000100", "10110111" ),
        ( "000011111", "10111101", "11010001" ),
        ( "011110001", "11011011", "11010101" ),
        ( "000001000", "10100000", "11101010" ),
        ( "011111100", "11110111", "11010101" ),
        ( "010011000", "11010111", "11101110" ),
        ( "001111000", "11101010", "11110110" ),
        ( "010110001", "01100111", "11110110" ),
        ( "011010010", "00111011", "10100011" ),
        ( "011110000", "10011111", "01111011" ),
        ( "001000100", "10011111", "00101000" ),
        ( "101001011", "11001100", "10110100" ),
        ( "100010111", "10010101", "11110011" ),
        ( "001001111", "11100100", "11001010" ),
        ( "100011101", "10000001", "11101111" ),
        ( "100000011", "01011000", "10011111" ),
        ( "101100000", "01011111", "11100011" ),
        ( "100110100", "11011010", "11111111" ),
        ( "001011100", "11010011", "11011111" ),
        ( "001101001", "11011000", "10100100" ),
        ( "100110100", "01111101", "10101011" ),
        ( "000110001", "11110101", "10001000" ),
        ( "000111000", "11100000", "11000111" ),
        ( "100001001", "11000111", "11110011" ),
        ( "101100100", "11000101", "00111010" ),
        ( "010011111", "10101110", "11011011" ),
        ( "001100001", "11010101", "00011111" ),
        ( "011110000", "10111110", "11110011" ),
        ( "010110100", "01001000", "11111010" ),
        ( "010101000", "11001110", "11101111" ),
        ( "001101011", "01110101", "01101000" ),
        ( "011110100", "11000100", "11100010" ),
        ( "011000100", "11001111", "11001011" ),
        ( "010001111", "01110001", "01010001" ),
        ( "101010011", "11010100", "11101111" ),
        ( "000100110", "11001111", "11111001" ),
        ( "100100011", "10111101", "11010001" ),
        ( "011100001", "01010001", "11001111" ),
        ( "100101000", "10010010", "10001000" ),
        ( "011110110", "01100111", "11000011" ),
        ( "001101001", "11100111", "01100000" ),
        ( "011011111", "01100111", "11011110" ),
        ( "101001111", "11011101", "11100111" ),
        ( "001000000", "11001011", "10111000" ),
        ( "000101000", "00101100", "00110100" ),
        ( "001110000", "11111100", "10101110" ),
        ( "010001010", "10011010", "10011000" ),
        ( "100100101", "00011111", "11010001" ),
        ( "100101010", "10010110", "11110111" ),
        ( "001011100", "11010110", "01101100" ),
        ( "000100001", "11111101", "11110100" ),
        ( "011010011", "11010001", "11010110" ),
        ( "010011000", "00111111", "11011010" ),
        ( "010001111", "11000111", "10100100" ),
        ( "011110011", "11101000", "10001010" ),
        ( "010100010", "11101111", "11110000" ),
        ( "001100011", "01000110", "01010000" ),
        ( "000011100", "11100100", "11101011" ),
        ( "001000010", "10011111", "11010100" ),
        ( "011111010", "10101101", "01100001" ),
        ( "011001010", "10110001", "10000001" ),
        ( "001101011", "10101101", "11011001" ),
        ( "001110010", "11100100", "11000100" ),
        ( "100101100", "00010100", "11011100" ),
        ( "000100100", "10010101", "11111110" ),
        ( "100001101", "11000111", "01111100" ),
        ( "010001010", "10100111", "11001111" ),
        ( "011011110", "11101101", "10001110" ),
        ( "000101111", "11110011", "11101010" ),
        ( "001100110", "10110111", "11111001" ),
        ( "100101110", "11011011", "10000011" ),
        ( "011011111", "10110001", "01000101" ),
        ( "000110011", "01101000", "11110010" ),
        ( "000111001", "00111101", "10110111" ),
        ( "011100101", "11110001", "11001010" ),
        ( "011000000", "10101000", "01000111" ),
        ( "101100000", "11001110", "10101111" ),
        ( "001101001", "01010011", "10000100" ),
        ( "001011010", "10000111", "11101011" ),
        ( "011010001", "01110101", "10110010" ),
        ( "010100001", "10111110", "11100000" ),
        ( "100011111", "10110001", "11010101" ),
        ( "101000011", "11110010", "11100010" ),
        ( "001011001", "10011100", "00111110" ),
        ( "010101111", "01110100", "10010000" ),
        ( "011001100", "11111001", "10000001" ),
        ( "001101111", "11011101", "01101010" ),
        ( "001001110", "10010010", "11001000" ),
        ( "000010100", "10111101", "11000011" ),
        ( "010100001", "01111101", "11001110" ),
        ( "010010100", "00101101", "01011111" ),
        ( "011110000", "11010001", "10110100" ),
        ( "011100111", "11000001", "11000111" ),
        ( "101001111", "11111011", "10100001" ),
        ( "100110111", "10010110", "10111011" ),
        ( "000001100", "10001011", "10010010" ),
        ( "101000110", "11010100", "11010110" ),
        ( "010011111", "11100010", "11111111" ),
        ( "010101011", "11111011", "10001010" )
    );

    constant check_result : boolean := true;

    component rgb2hsv is
        port(
            clk        : in  STD_LOGIC;
            rstn       : in  STD_LOGIC;
            data_rdy   : in  STD_LOGIC;
            r          : in  STD_LOGIC_VECTOR(7 downto 0);
            g          : in  STD_LOGIC_VECTOR(7 downto 0);
            b          : in  STD_LOGIC_VECTOR(7 downto 0);
            result_rdy : out STD_LOGIC;
            h          : out STD_LOGIC_VECTOR(8 downto 0);
            s          : out STD_LOGIC_VECTOR(7 downto 0);
            v          : out STD_LOGIC_VECTOR(7 downto 0)
        );
    end component;

    signal clk        : STD_LOGIC  := '1';
    signal rstn       : STD_LOGIC;
    signal data_rdy   : STD_LOGIC;
    signal r          : STD_LOGIC_VECTOR(7 downto 0);
    signal g          : STD_LOGIC_VECTOR(7 downto 0);
    signal b          : STD_LOGIC_VECTOR(7 downto 0);
    signal result_rdy : STD_LOGIC;
    signal h          : STD_LOGIC_VECTOR(8 downto 0);
    signal s          : STD_LOGIC_VECTOR(7 downto 0);
    signal v          : STD_LOGIC_VECTOR(7 downto 0);

begin

    UUT : rgb2hsv
        port map(
            clk        => clk,
            rstn       => rstn,
            data_rdy   => data_rdy,
            r          => r,
            g          => g,
            b          => b,
            result_rdy => result_rdy,
            h          => h,
            s          => s,
            v          => v
        );


    STIMULI_GEN : process
    begin

        rstn     <= '0';
        data_rdy <= '0';
        r        <= X"00";
        g        <= X"00";
        b        <= X"00";

        wait for 100 ns;
        wait until falling_edge(clk);

        rstn     <= '1';
        wait until falling_edge(clk);
    
        input_start <= cycle_counter;
        for i in 0 to 50 loop
            r        <= rgb_data(i).r;
            g        <= rgb_data(i).g;
            b        <= rgb_data(i).b;
            data_rdy <= '1';
            wait until falling_edge(clk);
        end loop;

        --
        data_rdy <= '0';
        wait until falling_edge(clk);
        wait until falling_edge(clk);
        wait until falling_edge(clk);
        wait until falling_edge(clk);
        wait until falling_edge(clk);

        for i in 51 to rgb_data'length-1 loop
            r        <= rgb_data(i).r;
            g        <= rgb_data(i).g;
            b        <= rgb_data(i).b;
            data_rdy <= '1';
            wait until falling_edge(clk);
        end loop;
        data_rdy <= '0';
        wait;
    end process;

    RESULT_TEST : process
    begin
        if check_result then
            if rstn /= '1' then
                wait until rstn = '1';
            end if;
            index <= 0;
            while index < hsv_data'length loop
                wait until falling_edge(clk);
                if result_rdy = '1' then
            if index = 0 then
            output_start <= cycle_counter;
            end if;

                    assert
                        (h = hsv_data(index).h) and (s = hsv_data(index).s) and (v = hsv_data(index).v)
                        report "error in hsv data - "
                            & "index: " & integer'image(index)
                            & "r: " & integer'image(conv_integer(rgb_data(index).r))
                            & ", g: " & integer'image(conv_integer(rgb_data(index).g))
                            & ", b: " & integer'image(conv_integer(rgb_data(index).b))
                            & ", h: " & integer'image(conv_integer(h)) & " ?= "  & integer'image(conv_integer(hsv_data(index).h))
                            & ", s: " & integer'image(conv_integer(s)) & " ?= "  & integer'image(conv_integer(hsv_data(index).s))
                            & ", v: " & integer'image(conv_integer(v)) & " ?= "  & integer'image(conv_integer(hsv_data(index).v))
                        severity failure;
                    index <= index + 1;
                end if;
            end loop;
            assert true report "all data correct" severity note;
            while true loop
                wait until falling_edge(clk);
                if result_rdy = '1' then
                    assert false report "extra result received" severity error;
                end if;
            end loop;
        end if;
        wait;
    end process;


    check_result_count: process
    begin        
        wait for 12100 ns; 
                
        assert index >= hsv_data'length
                report "Component did not generate the expected number of results!"
                severity failure;
        
        report "The pipeline length of the component is: " & integer'image(output_start - input_start);

        assert (output_start - input_start) >= 10
                report "Component is not pipelined properly!"
                severity failure;
                
        
        report "Test sucessful!";
        
        wait;
    end process;


    CLK_GEN : process(clk)
    begin
        clk <= not clk after 5 ns;
    if clk = '1' then
        cycle_counter <= cycle_counter + 1;
    end if;
    end process;

end architecture rtl;
